library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity scan is
   port (
      -- Clock
      clk_i      : in  std_logic;

      scan_i     : in  std_logic_vector(7 downto 0);
      ascii_o    : out std_logic_vector(7 downto 0)
   );
end scan;

architecture Structural of scan is

   type t_rom is array (0 to 255) of std_logic_vector(7 downto 0);

   constant scancode_rom : t_rom := (
      X"00",   -- 00
      X"00",   -- 01
      X"00",   -- 02
      X"00",   -- 03
      X"00",   -- 04
      X"00",   -- 05
      X"00",   -- 06
      X"00",   -- 07
      X"00",   -- 08
      X"00",   -- 09
      X"00",   -- 0A
      X"00",   -- 0B
      X"00",   -- 0C
      X"00",   -- 0D
      X"00",   -- 0E
      X"00",   -- 0F

      X"00",   -- 10
      X"00",   -- 11
      X"00",   -- 12
      X"00",   -- 13
      X"00",   -- 14
      X"51",   -- 15
      X"31",   -- 16
      X"00",   -- 17
      X"00",   -- 18
      X"00",   -- 19
      X"5A",   -- 1A
      X"53",   -- 1B
      X"41",   -- 1C
      X"57",   -- 1D
      X"32",   -- 1E
      X"00",   -- 1F

      X"00",   -- 20
      X"43",   -- 21
      X"58",   -- 22
      X"44",   -- 23
      X"45",   -- 24
      X"34",   -- 25
      X"33",   -- 26
      X"00",   -- 27
      X"00",   -- 28
      X"20",   -- 29
      X"56",   -- 2A
      X"46",   -- 2B
      X"54",   -- 2C
      X"52",   -- 2D
      X"35",   -- 2E
      X"00",   -- 2F

      X"00",   -- 30
      X"4E",   -- 31
      X"42",   -- 32
      X"48",   -- 33
      X"47",   -- 34
      X"59",   -- 35
      X"36",   -- 36
      X"00",   -- 37
      X"00",   -- 38
      X"00",   -- 39
      X"4D",   -- 3A
      X"4A",   -- 3B
      X"55",   -- 3C
      X"37",   -- 3D
      X"38",   -- 3E
      X"00",   -- 3F

      X"00",   -- 40
      X"00",   -- 41
      X"4B",   -- 42
      X"49",   -- 43
      X"4F",   -- 44
      X"30",   -- 45
      X"39",   -- 46
      X"00",   -- 47
      X"00",   -- 48
      X"00",   -- 49
      X"00",   -- 4A
      X"4C",   -- 4B
      X"00",   -- 4C
      X"50",   -- 4D
      X"00",   -- 4E
      X"00",   -- 4F

      X"00",   -- 50
      X"00",   -- 51
      X"00",   -- 52
      X"00",   -- 53
      X"00",   -- 54
      X"00",   -- 55
      X"00",   -- 56
      X"00",   -- 57
      X"00",   -- 58
      X"00",   -- 59
      X"00",   -- 5A
      X"00",   -- 5B
      X"00",   -- 5C
      X"00",   -- 5D
      X"00",   -- 5E
      X"00",   -- 5F

      X"00",   -- 60
      X"00",   -- 61
      X"00",   -- 62
      X"00",   -- 63
      X"00",   -- 64
      X"00",   -- 65
      X"00",   -- 66
      X"00",   -- 67
      X"00",   -- 68
      X"00",   -- 69
      X"00",   -- 6A
      X"00",   -- 6B
      X"00",   -- 6C
      X"00",   -- 6D
      X"00",   -- 6E
      X"00",   -- 6F

      X"00",   -- 70
      X"00",   -- 71
      X"00",   -- 72
      X"00",   -- 73
      X"00",   -- 74
      X"00",   -- 75
      X"00",   -- 76
      X"00",   -- 77
      X"00",   -- 78
      X"00",   -- 79
      X"00",   -- 7A
      X"00",   -- 7B
      X"00",   -- 7C
      X"00",   -- 7D
      X"00",   -- 7E
      X"00",   -- 7F

      X"00",   -- 80
      X"00",   -- 81
      X"00",   -- 82
      X"00",   -- 83
      X"00",   -- 84
      X"00",   -- 85
      X"00",   -- 86
      X"00",   -- 87
      X"00",   -- 88
      X"00",   -- 89
      X"00",   -- 8A
      X"00",   -- 8B
      X"00",   -- 8C
      X"00",   -- 8D
      X"00",   -- 8E
      X"00",   -- 8F

      X"00",   -- 90
      X"00",   -- 91
      X"00",   -- 92
      X"00",   -- 93
      X"00",   -- 94
      X"00",   -- 95
      X"00",   -- 96
      X"00",   -- 97
      X"00",   -- 98
      X"00",   -- 99
      X"00",   -- 9A
      X"00",   -- 9B
      X"00",   -- 9C
      X"00",   -- 9D
      X"00",   -- 9E
      X"00",   -- 9F

      X"00",   -- A0
      X"00",   -- A1
      X"00",   -- A2
      X"00",   -- A3
      X"00",   -- A4
      X"00",   -- A5
      X"00",   -- A6
      X"00",   -- A7
      X"00",   -- A8
      X"00",   -- A9
      X"00",   -- AA
      X"00",   -- AB
      X"00",   -- AC
      X"00",   -- AD
      X"00",   -- AE
      X"00",   -- AF

      X"00",   -- B0
      X"00",   -- B1
      X"00",   -- B2
      X"00",   -- B3
      X"00",   -- B4
      X"00",   -- B5
      X"00",   -- B6
      X"00",   -- B7
      X"00",   -- B8
      X"00",   -- B9
      X"00",   -- BA
      X"00",   -- BB
      X"00",   -- BC
      X"00",   -- BD
      X"00",   -- BE
      X"00",   -- BF

      X"00",   -- C0
      X"00",   -- C1
      X"00",   -- C2
      X"00",   -- C3
      X"00",   -- C4
      X"00",   -- C5
      X"00",   -- C6
      X"00",   -- C7
      X"00",   -- C8
      X"00",   -- C9
      X"00",   -- CA
      X"00",   -- CB
      X"00",   -- CC
      X"00",   -- CD
      X"00",   -- CE
      X"00",   -- CF

      X"00",   -- D0
      X"00",   -- D1
      X"00",   -- D2
      X"00",   -- D3
      X"00",   -- D4
      X"00",   -- D5
      X"00",   -- D6
      X"00",   -- D7
      X"00",   -- D8
      X"00",   -- D9
      X"00",   -- DA
      X"00",   -- DB
      X"00",   -- DC
      X"00",   -- DD
      X"00",   -- DE
      X"00",   -- DF

      X"00",   -- E0
      X"00",   -- E1
      X"00",   -- E2
      X"00",   -- E3
      X"00",   -- E4
      X"00",   -- E5
      X"00",   -- E6
      X"00",   -- E7
      X"00",   -- E8
      X"00",   -- E9
      X"00",   -- EA
      X"00",   -- EB
      X"00",   -- EC
      X"00",   -- ED
      X"00",   -- EE
      X"00",   -- EF

      X"00",   -- F0
      X"00",   -- F1
      X"00",   -- F2
      X"00",   -- F3
      X"00",   -- F4
      X"00",   -- F5
      X"00",   -- F6
      X"00",   -- F7
      X"00",   -- F8
      X"00",   -- F9
      X"00",   -- FA
      X"00",   -- FB
      X"00",   -- FC
      X"00",   -- FD
      X"00",   -- FE
      X"00"    -- FF
   );

begin

end Structural;


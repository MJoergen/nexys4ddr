library ieee;
use ieee.std_logic_1164.all;

-- Eventually, this block will handle the interface between the CPU and the
-- VERA, i.e. translate the CPU memory map into reads and writes to the VERA.
--
-- But for now, since there is no CPU, this block has a list of hardcoded
-- writes that it executes once at startup. These writes are gathered by
-- running the x16-emulator and having it dump all the writes to VERA.  There
-- were additional writes to clear the screen, but I've left them out, in order
-- to keep this file to a manageable size. Instead, I've simulated the clearing
-- of the screen by intializing the entire Video RAM to the value 0x66, which
-- corresponds to the blue colour, see vram.vhd.

entity cpu is
   port (
      clk_i     : in  std_logic;

      -- These will be connected to the vram block.
      -- TBD: What about the configuration settings, i.e. 0xFxxxx?
      wr_addr_o : out std_logic_vector(16 downto 0);
      wr_en_o   : out std_logic;
      wr_data_o : out std_logic_vector( 7 downto 0)
   );
end cpu;

architecture structural of cpu is

   -- This defines a type containing an array of bytes
   type wr_record is record
      addr : std_logic_vector(15 downto 0);
      data : std_logic_vector( 7 downto 0);
   end record wr_record;
   type wr_record_vector is array (natural range <>) of wr_record;

   constant wr_default : wr_record_vector := (
      -- The first part is the map area, i.e. the characters and colours.
      (X"0000", X"5F"),
      (X"0001", X"64"),
      (X"0002", X"A0"),
      (X"0003", X"64"),
      (X"0004", X"A0"),
      (X"0005", X"64"),
      (X"0006", X"DF"),
      (X"0007", X"64"),
      (X"0008", X"20"),
      (X"0009", X"64"),
      (X"000A", X"20"),
      (X"000B", X"64"),
      (X"000C", X"20"),
      (X"000D", X"64"),
      (X"000E", X"E9"),
      (X"000F", X"64"),
      (X"0010", X"A0"),
      (X"0011", X"64"),
      (X"0012", X"A0"),
      (X"0013", X"64"),
      (X"0014", X"69"),
      (X"0015", X"64"),
      (X"0100", X"20"),
      (X"0101", X"6E"),
      (X"0102", X"5F"),
      (X"0103", X"6E"),
      (X"0104", X"A0"),
      (X"0105", X"6E"),
      (X"0106", X"A0"),
      (X"0107", X"6E"),
      (X"0108", X"DF"),
      (X"0109", X"6E"),
      (X"010A", X"20"),
      (X"010B", X"6E"),
      (X"010C", X"E9"),
      (X"010D", X"6E"),
      (X"010E", X"A0"),
      (X"010F", X"6E"),
      (X"0110", X"A0"),
      (X"0111", X"6E"),
      (X"0112", X"69"),
      (X"0113", X"6E"),
      (X"0114", X"20"),
      (X"0115", X"61"),
      (X"0116", X"20"),
      (X"0117", X"61"),
      (X"0118", X"2A"),
      (X"0119", X"61"),
      (X"011A", X"2A"),
      (X"011B", X"61"),
      (X"011C", X"2A"),
      (X"011D", X"61"),
      (X"011E", X"2A"),
      (X"011F", X"61"),
      (X"0120", X"20"),
      (X"0121", X"61"),
      (X"0122", X"03"),
      (X"0123", X"61"),
      (X"0124", X"0F"),
      (X"0125", X"61"),
      (X"0126", X"0D"),
      (X"0127", X"61"),
      (X"0128", X"0D"),
      (X"0129", X"61"),
      (X"012A", X"01"),
      (X"012B", X"61"),
      (X"012C", X"0E"),
      (X"012D", X"61"),
      (X"012E", X"04"),
      (X"012F", X"61"),
      (X"0130", X"05"),
      (X"0131", X"61"),
      (X"0132", X"12"),
      (X"0133", X"61"),
      (X"0134", X"20"),
      (X"0135", X"61"),
      (X"0136", X"18"),
      (X"0137", X"61"),
      (X"0138", X"31"),
      (X"0139", X"61"),
      (X"013A", X"36"),
      (X"013B", X"61"),
      (X"013C", X"20"),
      (X"013D", X"61"),
      (X"013E", X"02"),
      (X"013F", X"61"),
      (X"0140", X"01"),
      (X"0141", X"61"),
      (X"0142", X"13"),
      (X"0143", X"61"),
      (X"0144", X"09"),
      (X"0145", X"61"),
      (X"0146", X"03"),
      (X"0147", X"61"),
      (X"0148", X"20"),
      (X"0149", X"61"),
      (X"014A", X"16"),
      (X"014B", X"61"),
      (X"014C", X"32"),
      (X"014D", X"61"),
      (X"014E", X"20"),
      (X"014F", X"61"),
      (X"0150", X"2A"),
      (X"0151", X"61"),
      (X"0152", X"2A"),
      (X"0153", X"61"),
      (X"0154", X"2A"),
      (X"0155", X"61"),
      (X"0156", X"2A"),
      (X"0157", X"61"),
      (X"0200", X"20"),
      (X"0201", X"63"),
      (X"0202", X"20"),
      (X"0203", X"63"),
      (X"0204", X"5F"),
      (X"0205", X"63"),
      (X"0206", X"A0"),
      (X"0207", X"63"),
      (X"0208", X"A0"),
      (X"0209", X"63"),
      (X"020A", X"20"),
      (X"020B", X"63"),
      (X"020C", X"A0"),
      (X"020D", X"63"),
      (X"020E", X"A0"),
      (X"020F", X"63"),
      (X"0210", X"69"),
      (X"0211", X"63"),
      (X"0300", X"20"),
      (X"0301", X"65"),
      (X"0302", X"20"),
      (X"0303", X"65"),
      (X"0304", X"20"),
      (X"0305", X"65"),
      (X"0306", X"20"),
      (X"0307", X"65"),
      (X"0308", X"A0"),
      (X"0309", X"65"),
      (X"030A", X"20"),
      (X"030B", X"65"),
      (X"030C", X"A0"),
      (X"030D", X"65"),
      (X"030E", X"20"),
      (X"030F", X"61"),
      (X"0310", X"20"),
      (X"0311", X"61"),
      (X"0312", X"20"),
      (X"0313", X"61"),
      (X"0314", X"20"),
      (X"0315", X"61"),
      (X"0316", X"20"),
      (X"0317", X"61"),
      (X"0318", X"35"),
      (X"0319", X"61"),
      (X"031A", X"31"),
      (X"031B", X"61"),
      (X"031C", X"32"),
      (X"031D", X"61"),
      (X"031E", X"0B"),
      (X"031F", X"61"),
      (X"0320", X"20"),
      (X"0321", X"61"),
      (X"0322", X"08"),
      (X"0323", X"61"),
      (X"0324", X"09"),
      (X"0325", X"61"),
      (X"0326", X"07"),
      (X"0327", X"61"),
      (X"0328", X"08"),
      (X"0329", X"61"),
      (X"032A", X"20"),
      (X"032B", X"61"),
      (X"032C", X"12"),
      (X"032D", X"61"),
      (X"032E", X"01"),
      (X"032F", X"61"),
      (X"0330", X"0D"),
      (X"0331", X"61"),
      (X"0400", X"20"),
      (X"0401", X"67"),
      (X"0402", X"20"),
      (X"0403", X"67"),
      (X"0404", X"E9"),
      (X"0405", X"67"),
      (X"0406", X"A0"),
      (X"0407", X"67"),
      (X"0408", X"A0"),
      (X"0409", X"67"),
      (X"040A", X"20"),
      (X"040B", X"67"),
      (X"040C", X"A0"),
      (X"040D", X"67"),
      (X"040E", X"A0"),
      (X"040F", X"67"),
      (X"0410", X"DF"),
      (X"0411", X"67"),
      (X"0500", X"20"),
      (X"0501", X"68"),
      (X"0502", X"E9"),
      (X"0503", X"68"),
      (X"0504", X"A0"),
      (X"0505", X"68"),
      (X"0506", X"A0"),
      (X"0507", X"68"),
      (X"0508", X"69"),
      (X"0509", X"68"),
      (X"050A", X"20"),
      (X"050B", X"68"),
      (X"050C", X"5F"),
      (X"050D", X"68"),
      (X"050E", X"A0"),
      (X"050F", X"68"),
      (X"0510", X"A0"),
      (X"0511", X"68"),
      (X"0512", X"DF"),
      (X"0513", X"68"),
      (X"0514", X"20"),
      (X"0515", X"61"),
      (X"0516", X"20"),
      (X"0517", X"61"),
      (X"0518", X"33"),
      (X"0519", X"61"),
      (X"051A", X"38"),
      (X"051B", X"61"),
      (X"051C", X"36"),
      (X"051D", X"61"),
      (X"051E", X"35"),
      (X"051F", X"61"),
      (X"0520", X"35"),
      (X"0521", X"61"),
      (X"0522", X"20"),
      (X"0523", X"61"),
      (X"0524", X"02"),
      (X"0525", X"61"),
      (X"0526", X"01"),
      (X"0527", X"61"),
      (X"0528", X"13"),
      (X"0529", X"61"),
      (X"052A", X"09"),
      (X"052B", X"61"),
      (X"052C", X"03"),
      (X"052D", X"61"),
      (X"052E", X"20"),
      (X"052F", X"61"),
      (X"0530", X"02"),
      (X"0531", X"61"),
      (X"0532", X"19"),
      (X"0533", X"61"),
      (X"0534", X"14"),
      (X"0535", X"61"),
      (X"0536", X"05"),
      (X"0537", X"61"),
      (X"0538", X"13"),
      (X"0539", X"61"),
      (X"053A", X"20"),
      (X"053B", X"61"),
      (X"053C", X"06"),
      (X"053D", X"61"),
      (X"053E", X"12"),
      (X"053F", X"61"),
      (X"0540", X"05"),
      (X"0541", X"61"),
      (X"0542", X"05"),
      (X"0543", X"61"),
      (X"0600", X"E9"),
      (X"0601", X"62"),
      (X"0602", X"A0"),
      (X"0603", X"62"),
      (X"0604", X"A0"),
      (X"0605", X"62"),
      (X"0606", X"69"),
      (X"0607", X"62"),
      (X"0608", X"20"),
      (X"0609", X"62"),
      (X"060A", X"20"),
      (X"060B", X"62"),
      (X"060C", X"20"),
      (X"060D", X"62"),
      (X"060E", X"5F"),
      (X"060F", X"62"),
      (X"0610", X"A0"),
      (X"0611", X"62"),
      (X"0612", X"A0"),
      (X"0613", X"62"),
      (X"0614", X"DF"),
      (X"0615", X"62"),
      (X"0800", X"12"),
      (X"0801", X"61"),
      (X"0802", X"05"),
      (X"0803", X"61"),
      (X"0804", X"01"),
      (X"0805", X"61"),
      (X"0806", X"04"),
      (X"0807", X"61"),
      (X"0808", X"19"),
      (X"0809", X"61"),
      (X"080A", X"2E"),
      (X"080B", X"61"),

      -- The second part is the tile map, i.e. the font
      (X"F800", X"3C"),
      (X"F801", X"66"),
      (X"F802", X"6E"),
      (X"F803", X"6E"),
      (X"F804", X"60"),
      (X"F805", X"62"),
      (X"F806", X"3C"),
      (X"F807", X"00"),
      (X"F808", X"18"),
      (X"F809", X"3C"),
      (X"F80A", X"66"),
      (X"F80B", X"7E"),
      (X"F80C", X"66"),
      (X"F80D", X"66"),
      (X"F80E", X"66"),
      (X"F80F", X"00"),
      (X"F810", X"7C"),
      (X"F811", X"66"),
      (X"F812", X"66"),
      (X"F813", X"7C"),
      (X"F814", X"66"),
      (X"F815", X"66"),
      (X"F816", X"7C"),
      (X"F817", X"00"),
      (X"F818", X"3C"),
      (X"F819", X"66"),
      (X"F81A", X"60"),
      (X"F81B", X"60"),
      (X"F81C", X"60"),
      (X"F81D", X"66"),
      (X"F81E", X"3C"),
      (X"F81F", X"00"),
      (X"F820", X"78"),
      (X"F821", X"6C"),
      (X"F822", X"66"),
      (X"F823", X"66"),
      (X"F824", X"66"),
      (X"F825", X"6C"),
      (X"F826", X"78"),
      (X"F827", X"00"),
      (X"F828", X"7E"),
      (X"F829", X"60"),
      (X"F82A", X"60"),
      (X"F82B", X"78"),
      (X"F82C", X"60"),
      (X"F82D", X"60"),
      (X"F82E", X"7E"),
      (X"F82F", X"00"),
      (X"F830", X"7E"),
      (X"F831", X"60"),
      (X"F832", X"60"),
      (X"F833", X"78"),
      (X"F834", X"60"),
      (X"F835", X"60"),
      (X"F836", X"60"),
      (X"F837", X"00"),
      (X"F838", X"3C"),
      (X"F839", X"66"),
      (X"F83A", X"60"),
      (X"F83B", X"6E"),
      (X"F83C", X"66"),
      (X"F83D", X"66"),
      (X"F83E", X"3C"),
      (X"F83F", X"00"),
      (X"F840", X"66"),
      (X"F841", X"66"),
      (X"F842", X"66"),
      (X"F843", X"7E"),
      (X"F844", X"66"),
      (X"F845", X"66"),
      (X"F846", X"66"),
      (X"F847", X"00"),
      (X"F848", X"3C"),
      (X"F849", X"18"),
      (X"F84A", X"18"),
      (X"F84B", X"18"),
      (X"F84C", X"18"),
      (X"F84D", X"18"),
      (X"F84E", X"3C"),
      (X"F84F", X"00"),
      (X"F850", X"1E"),
      (X"F851", X"0C"),
      (X"F852", X"0C"),
      (X"F853", X"0C"),
      (X"F854", X"0C"),
      (X"F855", X"6C"),
      (X"F856", X"38"),
      (X"F857", X"00"),
      (X"F858", X"66"),
      (X"F859", X"6C"),
      (X"F85A", X"78"),
      (X"F85B", X"70"),
      (X"F85C", X"78"),
      (X"F85D", X"6C"),
      (X"F85E", X"66"),
      (X"F85F", X"00"),
      (X"F860", X"60"),
      (X"F861", X"60"),
      (X"F862", X"60"),
      (X"F863", X"60"),
      (X"F864", X"60"),
      (X"F865", X"60"),
      (X"F866", X"7E"),
      (X"F867", X"00"),
      (X"F868", X"63"),
      (X"F869", X"77"),
      (X"F86A", X"7F"),
      (X"F86B", X"6B"),
      (X"F86C", X"63"),
      (X"F86D", X"63"),
      (X"F86E", X"63"),
      (X"F86F", X"00"),
      (X"F870", X"66"),
      (X"F871", X"76"),
      (X"F872", X"7E"),
      (X"F873", X"7E"),
      (X"F874", X"6E"),
      (X"F875", X"66"),
      (X"F876", X"66"),
      (X"F877", X"00"),
      (X"F878", X"3C"),
      (X"F879", X"66"),
      (X"F87A", X"66"),
      (X"F87B", X"66"),
      (X"F87C", X"66"),
      (X"F87D", X"66"),
      (X"F87E", X"3C"),
      (X"F87F", X"00"),
      (X"F880", X"7C"),
      (X"F881", X"66"),
      (X"F882", X"66"),
      (X"F883", X"7C"),
      (X"F884", X"60"),
      (X"F885", X"60"),
      (X"F886", X"60"),
      (X"F887", X"00"),
      (X"F888", X"3C"),
      (X"F889", X"66"),
      (X"F88A", X"66"),
      (X"F88B", X"66"),
      (X"F88C", X"66"),
      (X"F88D", X"3C"),
      (X"F88E", X"0E"),
      (X"F88F", X"00"),
      (X"F890", X"7C"),
      (X"F891", X"66"),
      (X"F892", X"66"),
      (X"F893", X"7C"),
      (X"F894", X"78"),
      (X"F895", X"6C"),
      (X"F896", X"66"),
      (X"F897", X"00"),
      (X"F898", X"3C"),
      (X"F899", X"66"),
      (X"F89A", X"60"),
      (X"F89B", X"3C"),
      (X"F89C", X"06"),
      (X"F89D", X"66"),
      (X"F89E", X"3C"),
      (X"F89F", X"00"),
      (X"F8A0", X"7E"),
      (X"F8A1", X"18"),
      (X"F8A2", X"18"),
      (X"F8A3", X"18"),
      (X"F8A4", X"18"),
      (X"F8A5", X"18"),
      (X"F8A6", X"18"),
      (X"F8A7", X"00"),
      (X"F8A8", X"66"),
      (X"F8A9", X"66"),
      (X"F8AA", X"66"),
      (X"F8AB", X"66"),
      (X"F8AC", X"66"),
      (X"F8AD", X"66"),
      (X"F8AE", X"3C"),
      (X"F8AF", X"00"),
      (X"F8B0", X"66"),
      (X"F8B1", X"66"),
      (X"F8B2", X"66"),
      (X"F8B3", X"66"),
      (X"F8B4", X"66"),
      (X"F8B5", X"3C"),
      (X"F8B6", X"18"),
      (X"F8B7", X"00"),
      (X"F8B8", X"63"),
      (X"F8B9", X"63"),
      (X"F8BA", X"63"),
      (X"F8BB", X"6B"),
      (X"F8BC", X"7F"),
      (X"F8BD", X"77"),
      (X"F8BE", X"63"),
      (X"F8BF", X"00"),
      (X"F8C0", X"66"),
      (X"F8C1", X"66"),
      (X"F8C2", X"3C"),
      (X"F8C3", X"18"),
      (X"F8C4", X"3C"),
      (X"F8C5", X"66"),
      (X"F8C6", X"66"),
      (X"F8C7", X"00"),
      (X"F8C8", X"66"),
      (X"F8C9", X"66"),
      (X"F8CA", X"66"),
      (X"F8CB", X"3C"),
      (X"F8CC", X"18"),
      (X"F8CD", X"18"),
      (X"F8CE", X"18"),
      (X"F8CF", X"00"),
      (X"F8D0", X"7E"),
      (X"F8D1", X"06"),
      (X"F8D2", X"0C"),
      (X"F8D3", X"18"),
      (X"F8D4", X"30"),
      (X"F8D5", X"60"),
      (X"F8D6", X"7E"),
      (X"F8D7", X"00"),
      (X"F8D8", X"3C"),
      (X"F8D9", X"30"),
      (X"F8DA", X"30"),
      (X"F8DB", X"30"),
      (X"F8DC", X"30"),
      (X"F8DD", X"30"),
      (X"F8DE", X"3C"),
      (X"F8DF", X"00"),
      (X"F8E0", X"0C"),
      (X"F8E1", X"12"),
      (X"F8E2", X"30"),
      (X"F8E3", X"7C"),
      (X"F8E4", X"30"),
      (X"F8E5", X"62"),
      (X"F8E6", X"FC"),
      (X"F8E7", X"00"),
      (X"F8E8", X"3C"),
      (X"F8E9", X"0C"),
      (X"F8EA", X"0C"),
      (X"F8EB", X"0C"),
      (X"F8EC", X"0C"),
      (X"F8ED", X"0C"),
      (X"F8EE", X"3C"),
      (X"F8EF", X"00"),
      (X"F8F0", X"00"),
      (X"F8F1", X"18"),
      (X"F8F2", X"3C"),
      (X"F8F3", X"7E"),
      (X"F8F4", X"18"),
      (X"F8F5", X"18"),
      (X"F8F6", X"18"),
      (X"F8F7", X"18"),
      (X"F8F8", X"00"),
      (X"F8F9", X"10"),
      (X"F8FA", X"30"),
      (X"F8FB", X"7F"),
      (X"F8FC", X"7F"),
      (X"F8FD", X"30"),
      (X"F8FE", X"10"),
      (X"F8FF", X"00"),
      (X"F900", X"00"),
      (X"F901", X"00"),
      (X"F902", X"00"),
      (X"F903", X"00"),
      (X"F904", X"00"),
      (X"F905", X"00"),
      (X"F906", X"00"),
      (X"F907", X"00"),
      (X"F908", X"18"),
      (X"F909", X"18"),
      (X"F90A", X"18"),
      (X"F90B", X"18"),
      (X"F90C", X"00"),
      (X"F90D", X"00"),
      (X"F90E", X"18"),
      (X"F90F", X"00"),
      (X"F910", X"66"),
      (X"F911", X"66"),
      (X"F912", X"66"),
      (X"F913", X"00"),
      (X"F914", X"00"),
      (X"F915", X"00"),
      (X"F916", X"00"),
      (X"F917", X"00"),
      (X"F918", X"66"),
      (X"F919", X"66"),
      (X"F91A", X"FF"),
      (X"F91B", X"66"),
      (X"F91C", X"FF"),
      (X"F91D", X"66"),
      (X"F91E", X"66"),
      (X"F91F", X"00"),
      (X"F920", X"18"),
      (X"F921", X"3E"),
      (X"F922", X"60"),
      (X"F923", X"3C"),
      (X"F924", X"06"),
      (X"F925", X"7C"),
      (X"F926", X"18"),
      (X"F927", X"00"),
      (X"F928", X"62"),
      (X"F929", X"66"),
      (X"F92A", X"0C"),
      (X"F92B", X"18"),
      (X"F92C", X"30"),
      (X"F92D", X"66"),
      (X"F92E", X"46"),
      (X"F92F", X"00"),
      (X"F930", X"3C"),
      (X"F931", X"66"),
      (X"F932", X"3C"),
      (X"F933", X"38"),
      (X"F934", X"67"),
      (X"F935", X"66"),
      (X"F936", X"3F"),
      (X"F937", X"00"),
      (X"F938", X"06"),
      (X"F939", X"0C"),
      (X"F93A", X"18"),
      (X"F93B", X"00"),
      (X"F93C", X"00"),
      (X"F93D", X"00"),
      (X"F93E", X"00"),
      (X"F93F", X"00"),
      (X"F940", X"0C"),
      (X"F941", X"18"),
      (X"F942", X"30"),
      (X"F943", X"30"),
      (X"F944", X"30"),
      (X"F945", X"18"),
      (X"F946", X"0C"),
      (X"F947", X"00"),
      (X"F948", X"30"),
      (X"F949", X"18"),
      (X"F94A", X"0C"),
      (X"F94B", X"0C"),
      (X"F94C", X"0C"),
      (X"F94D", X"18"),
      (X"F94E", X"30"),
      (X"F94F", X"00"),
      (X"F950", X"00"),
      (X"F951", X"66"),
      (X"F952", X"3C"),
      (X"F953", X"FF"),
      (X"F954", X"3C"),
      (X"F955", X"66"),
      (X"F956", X"00"),
      (X"F957", X"00"),
      (X"F958", X"00"),
      (X"F959", X"18"),
      (X"F95A", X"18"),
      (X"F95B", X"7E"),
      (X"F95C", X"18"),
      (X"F95D", X"18"),
      (X"F95E", X"00"),
      (X"F95F", X"00"),
      (X"F960", X"00"),
      (X"F961", X"00"),
      (X"F962", X"00"),
      (X"F963", X"00"),
      (X"F964", X"00"),
      (X"F965", X"18"),
      (X"F966", X"18"),
      (X"F967", X"30"),
      (X"F968", X"00"),
      (X"F969", X"00"),
      (X"F96A", X"00"),
      (X"F96B", X"7E"),
      (X"F96C", X"00"),
      (X"F96D", X"00"),
      (X"F96E", X"00"),
      (X"F96F", X"00"),
      (X"F970", X"00"),
      (X"F971", X"00"),
      (X"F972", X"00"),
      (X"F973", X"00"),
      (X"F974", X"00"),
      (X"F975", X"18"),
      (X"F976", X"18"),
      (X"F977", X"00"),
      (X"F978", X"00"),
      (X"F979", X"03"),
      (X"F97A", X"06"),
      (X"F97B", X"0C"),
      (X"F97C", X"18"),
      (X"F97D", X"30"),
      (X"F97E", X"60"),
      (X"F97F", X"00"),
      (X"F980", X"3C"),
      (X"F981", X"66"),
      (X"F982", X"6E"),
      (X"F983", X"76"),
      (X"F984", X"66"),
      (X"F985", X"66"),
      (X"F986", X"3C"),
      (X"F987", X"00"),
      (X"F988", X"18"),
      (X"F989", X"18"),
      (X"F98A", X"38"),
      (X"F98B", X"18"),
      (X"F98C", X"18"),
      (X"F98D", X"18"),
      (X"F98E", X"7E"),
      (X"F98F", X"00"),
      (X"F990", X"3C"),
      (X"F991", X"66"),
      (X"F992", X"06"),
      (X"F993", X"0C"),
      (X"F994", X"30"),
      (X"F995", X"60"),
      (X"F996", X"7E"),
      (X"F997", X"00"),
      (X"F998", X"3C"),
      (X"F999", X"66"),
      (X"F99A", X"06"),
      (X"F99B", X"1C"),
      (X"F99C", X"06"),
      (X"F99D", X"66"),
      (X"F99E", X"3C"),
      (X"F99F", X"00"),
      (X"F9A0", X"06"),
      (X"F9A1", X"0E"),
      (X"F9A2", X"1E"),
      (X"F9A3", X"66"),
      (X"F9A4", X"7F"),
      (X"F9A5", X"06"),
      (X"F9A6", X"06"),
      (X"F9A7", X"00"),
      (X"F9A8", X"7E"),
      (X"F9A9", X"60"),
      (X"F9AA", X"7C"),
      (X"F9AB", X"06"),
      (X"F9AC", X"06"),
      (X"F9AD", X"66"),
      (X"F9AE", X"3C"),
      (X"F9AF", X"00"),
      (X"F9B0", X"3C"),
      (X"F9B1", X"66"),
      (X"F9B2", X"60"),
      (X"F9B3", X"7C"),
      (X"F9B4", X"66"),
      (X"F9B5", X"66"),
      (X"F9B6", X"3C"),
      (X"F9B7", X"00"),
      (X"F9B8", X"7E"),
      (X"F9B9", X"66"),
      (X"F9BA", X"0C"),
      (X"F9BB", X"18"),
      (X"F9BC", X"18"),
      (X"F9BD", X"18"),
      (X"F9BE", X"18"),
      (X"F9BF", X"00"),
      (X"F9C0", X"3C"),
      (X"F9C1", X"66"),
      (X"F9C2", X"66"),
      (X"F9C3", X"3C"),
      (X"F9C4", X"66"),
      (X"F9C5", X"66"),
      (X"F9C6", X"3C"),
      (X"F9C7", X"00"),
      (X"F9C8", X"3C"),
      (X"F9C9", X"66"),
      (X"F9CA", X"66"),
      (X"F9CB", X"3E"),
      (X"F9CC", X"06"),
      (X"F9CD", X"66"),
      (X"F9CE", X"3C"),
      (X"F9CF", X"00"),
      (X"F9D0", X"00"),
      (X"F9D1", X"00"),
      (X"F9D2", X"18"),
      (X"F9D3", X"00"),
      (X"F9D4", X"00"),
      (X"F9D5", X"18"),
      (X"F9D6", X"00"),
      (X"F9D7", X"00"),
      (X"F9D8", X"00"),
      (X"F9D9", X"00"),
      (X"F9DA", X"18"),
      (X"F9DB", X"00"),
      (X"F9DC", X"00"),
      (X"F9DD", X"18"),
      (X"F9DE", X"18"),
      (X"F9DF", X"30"),
      (X"F9E0", X"0E"),
      (X"F9E1", X"18"),
      (X"F9E2", X"30"),
      (X"F9E3", X"60"),
      (X"F9E4", X"30"),
      (X"F9E5", X"18"),
      (X"F9E6", X"0E"),
      (X"F9E7", X"00"),
      (X"F9E8", X"00"),
      (X"F9E9", X"00"),
      (X"F9EA", X"7E"),
      (X"F9EB", X"00"),
      (X"F9EC", X"7E"),
      (X"F9ED", X"00"),
      (X"F9EE", X"00"),
      (X"F9EF", X"00"),
      (X"F9F0", X"70"),
      (X"F9F1", X"18"),
      (X"F9F2", X"0C"),
      (X"F9F3", X"06"),
      (X"F9F4", X"0C"),
      (X"F9F5", X"18"),
      (X"F9F6", X"70"),
      (X"F9F7", X"00"),
      (X"F9F8", X"3C"),
      (X"F9F9", X"66"),
      (X"F9FA", X"06"),
      (X"F9FB", X"0C"),
      (X"F9FC", X"18"),
      (X"F9FD", X"00"),
      (X"F9FE", X"18"),
      (X"F9FF", X"00"),
      (X"FA00", X"00"),
      (X"FA01", X"00"),
      (X"FA02", X"00"),
      (X"FA03", X"FF"),
      (X"FA04", X"FF"),
      (X"FA05", X"00"),
      (X"FA06", X"00"),
      (X"FA07", X"00"),
      (X"FA08", X"08"),
      (X"FA09", X"1C"),
      (X"FA0A", X"3E"),
      (X"FA0B", X"7F"),
      (X"FA0C", X"7F"),
      (X"FA0D", X"1C"),
      (X"FA0E", X"3E"),
      (X"FA0F", X"00"),
      (X"FA10", X"18"),
      (X"FA11", X"18"),
      (X"FA12", X"18"),
      (X"FA13", X"18"),
      (X"FA14", X"18"),
      (X"FA15", X"18"),
      (X"FA16", X"18"),
      (X"FA17", X"18"),
      (X"FA18", X"00"),
      (X"FA19", X"00"),
      (X"FA1A", X"00"),
      (X"FA1B", X"FF"),
      (X"FA1C", X"FF"),
      (X"FA1D", X"00"),
      (X"FA1E", X"00"),
      (X"FA1F", X"00"),
      (X"FA20", X"00"),
      (X"FA21", X"00"),
      (X"FA22", X"FF"),
      (X"FA23", X"FF"),
      (X"FA24", X"00"),
      (X"FA25", X"00"),
      (X"FA26", X"00"),
      (X"FA27", X"00"),
      (X"FA28", X"00"),
      (X"FA29", X"FF"),
      (X"FA2A", X"FF"),
      (X"FA2B", X"00"),
      (X"FA2C", X"00"),
      (X"FA2D", X"00"),
      (X"FA2E", X"00"),
      (X"FA2F", X"00"),
      (X"FA30", X"00"),
      (X"FA31", X"00"),
      (X"FA32", X"00"),
      (X"FA33", X"00"),
      (X"FA34", X"FF"),
      (X"FA35", X"FF"),
      (X"FA36", X"00"),
      (X"FA37", X"00"),
      (X"FA38", X"30"),
      (X"FA39", X"30"),
      (X"FA3A", X"30"),
      (X"FA3B", X"30"),
      (X"FA3C", X"30"),
      (X"FA3D", X"30"),
      (X"FA3E", X"30"),
      (X"FA3F", X"30"),
      (X"FA40", X"0C"),
      (X"FA41", X"0C"),
      (X"FA42", X"0C"),
      (X"FA43", X"0C"),
      (X"FA44", X"0C"),
      (X"FA45", X"0C"),
      (X"FA46", X"0C"),
      (X"FA47", X"0C"),
      (X"FA48", X"00"),
      (X"FA49", X"00"),
      (X"FA4A", X"00"),
      (X"FA4B", X"E0"),
      (X"FA4C", X"F0"),
      (X"FA4D", X"38"),
      (X"FA4E", X"18"),
      (X"FA4F", X"18"),
      (X"FA50", X"18"),
      (X"FA51", X"18"),
      (X"FA52", X"1C"),
      (X"FA53", X"0F"),
      (X"FA54", X"07"),
      (X"FA55", X"00"),
      (X"FA56", X"00"),
      (X"FA57", X"00"),
      (X"FA58", X"18"),
      (X"FA59", X"18"),
      (X"FA5A", X"38"),
      (X"FA5B", X"F0"),
      (X"FA5C", X"E0"),
      (X"FA5D", X"00"),
      (X"FA5E", X"00"),
      (X"FA5F", X"00"),
      (X"FA60", X"C0"),
      (X"FA61", X"C0"),
      (X"FA62", X"C0"),
      (X"FA63", X"C0"),
      (X"FA64", X"C0"),
      (X"FA65", X"C0"),
      (X"FA66", X"FF"),
      (X"FA67", X"FF"),
      (X"FA68", X"C0"),
      (X"FA69", X"E0"),
      (X"FA6A", X"70"),
      (X"FA6B", X"38"),
      (X"FA6C", X"1C"),
      (X"FA6D", X"0E"),
      (X"FA6E", X"07"),
      (X"FA6F", X"03"),
      (X"FA70", X"03"),
      (X"FA71", X"07"),
      (X"FA72", X"0E"),
      (X"FA73", X"1C"),
      (X"FA74", X"38"),
      (X"FA75", X"70"),
      (X"FA76", X"E0"),
      (X"FA77", X"C0"),
      (X"FA78", X"FF"),
      (X"FA79", X"FF"),
      (X"FA7A", X"C0"),
      (X"FA7B", X"C0"),
      (X"FA7C", X"C0"),
      (X"FA7D", X"C0"),
      (X"FA7E", X"C0"),
      (X"FA7F", X"C0"),
      (X"FA80", X"FF"),
      (X"FA81", X"FF"),
      (X"FA82", X"03"),
      (X"FA83", X"03"),
      (X"FA84", X"03"),
      (X"FA85", X"03"),
      (X"FA86", X"03"),
      (X"FA87", X"03"),
      (X"FA88", X"00"),
      (X"FA89", X"3C"),
      (X"FA8A", X"7E"),
      (X"FA8B", X"7E"),
      (X"FA8C", X"7E"),
      (X"FA8D", X"7E"),
      (X"FA8E", X"3C"),
      (X"FA8F", X"00"),
      (X"FA90", X"00"),
      (X"FA91", X"00"),
      (X"FA92", X"00"),
      (X"FA93", X"00"),
      (X"FA94", X"00"),
      (X"FA95", X"FF"),
      (X"FA96", X"FF"),
      (X"FA97", X"00"),
      (X"FA98", X"36"),
      (X"FA99", X"7F"),
      (X"FA9A", X"7F"),
      (X"FA9B", X"7F"),
      (X"FA9C", X"3E"),
      (X"FA9D", X"1C"),
      (X"FA9E", X"08"),
      (X"FA9F", X"00"),
      (X"FAA0", X"60"),
      (X"FAA1", X"60"),
      (X"FAA2", X"60"),
      (X"FAA3", X"60"),
      (X"FAA4", X"60"),
      (X"FAA5", X"60"),
      (X"FAA6", X"60"),
      (X"FAA7", X"60"),
      (X"FAA8", X"00"),
      (X"FAA9", X"00"),
      (X"FAAA", X"00"),
      (X"FAAB", X"07"),
      (X"FAAC", X"0F"),
      (X"FAAD", X"1C"),
      (X"FAAE", X"18"),
      (X"FAAF", X"18"),
      (X"FAB0", X"C3"),
      (X"FAB1", X"E7"),
      (X"FAB2", X"7E"),
      (X"FAB3", X"3C"),
      (X"FAB4", X"3C"),
      (X"FAB5", X"7E"),
      (X"FAB6", X"E7"),
      (X"FAB7", X"C3"),
      (X"FAB8", X"00"),
      (X"FAB9", X"3C"),
      (X"FABA", X"7E"),
      (X"FABB", X"66"),
      (X"FABC", X"66"),
      (X"FABD", X"7E"),
      (X"FABE", X"3C"),
      (X"FABF", X"00"),
      (X"FAC0", X"18"),
      (X"FAC1", X"18"),
      (X"FAC2", X"66"),
      (X"FAC3", X"66"),
      (X"FAC4", X"18"),
      (X"FAC5", X"18"),
      (X"FAC6", X"3C"),
      (X"FAC7", X"00"),
      (X"FAC8", X"06"),
      (X"FAC9", X"06"),
      (X"FACA", X"06"),
      (X"FACB", X"06"),
      (X"FACC", X"06"),
      (X"FACD", X"06"),
      (X"FACE", X"06"),
      (X"FACF", X"06"),
      (X"FAD0", X"08"),
      (X"FAD1", X"1C"),
      (X"FAD2", X"3E"),
      (X"FAD3", X"7F"),
      (X"FAD4", X"3E"),
      (X"FAD5", X"1C"),
      (X"FAD6", X"08"),
      (X"FAD7", X"00"),
      (X"FAD8", X"18"),
      (X"FAD9", X"18"),
      (X"FADA", X"18"),
      (X"FADB", X"FF"),
      (X"FADC", X"FF"),
      (X"FADD", X"18"),
      (X"FADE", X"18"),
      (X"FADF", X"18"),
      (X"FAE0", X"C0"),
      (X"FAE1", X"C0"),
      (X"FAE2", X"30"),
      (X"FAE3", X"30"),
      (X"FAE4", X"C0"),
      (X"FAE5", X"C0"),
      (X"FAE6", X"30"),
      (X"FAE7", X"30"),
      (X"FAE8", X"18"),
      (X"FAE9", X"18"),
      (X"FAEA", X"18"),
      (X"FAEB", X"18"),
      (X"FAEC", X"18"),
      (X"FAED", X"18"),
      (X"FAEE", X"18"),
      (X"FAEF", X"18"),
      (X"FAF0", X"00"),
      (X"FAF1", X"00"),
      (X"FAF2", X"03"),
      (X"FAF3", X"3E"),
      (X"FAF4", X"76"),
      (X"FAF5", X"36"),
      (X"FAF6", X"36"),
      (X"FAF7", X"00"),
      (X"FAF8", X"FF"),
      (X"FAF9", X"7F"),
      (X"FAFA", X"3F"),
      (X"FAFB", X"1F"),
      (X"FAFC", X"0F"),
      (X"FAFD", X"07"),
      (X"FAFE", X"03"),
      (X"FAFF", X"01"),
      (X"FB00", X"00"),
      (X"FB01", X"00"),
      (X"FB02", X"00"),
      (X"FB03", X"00"),
      (X"FB04", X"00"),
      (X"FB05", X"00"),
      (X"FB06", X"00"),
      (X"FB07", X"00"),
      (X"FB08", X"F0"),
      (X"FB09", X"F0"),
      (X"FB0A", X"F0"),
      (X"FB0B", X"F0"),
      (X"FB0C", X"F0"),
      (X"FB0D", X"F0"),
      (X"FB0E", X"F0"),
      (X"FB0F", X"F0"),
      (X"FB10", X"00"),
      (X"FB11", X"00"),
      (X"FB12", X"00"),
      (X"FB13", X"00"),
      (X"FB14", X"FF"),
      (X"FB15", X"FF"),
      (X"FB16", X"FF"),
      (X"FB17", X"FF"),
      (X"FB18", X"FF"),
      (X"FB19", X"00"),
      (X"FB1A", X"00"),
      (X"FB1B", X"00"),
      (X"FB1C", X"00"),
      (X"FB1D", X"00"),
      (X"FB1E", X"00"),
      (X"FB1F", X"00"),
      (X"FB20", X"00"),
      (X"FB21", X"00"),
      (X"FB22", X"00"),
      (X"FB23", X"00"),
      (X"FB24", X"00"),
      (X"FB25", X"00"),
      (X"FB26", X"00"),
      (X"FB27", X"FF"),
      (X"FB28", X"C0"),
      (X"FB29", X"C0"),
      (X"FB2A", X"C0"),
      (X"FB2B", X"C0"),
      (X"FB2C", X"C0"),
      (X"FB2D", X"C0"),
      (X"FB2E", X"C0"),
      (X"FB2F", X"C0"),
      (X"FB30", X"CC"),
      (X"FB31", X"CC"),
      (X"FB32", X"33"),
      (X"FB33", X"33"),
      (X"FB34", X"CC"),
      (X"FB35", X"CC"),
      (X"FB36", X"33"),
      (X"FB37", X"33"),
      (X"FB38", X"03"),
      (X"FB39", X"03"),
      (X"FB3A", X"03"),
      (X"FB3B", X"03"),
      (X"FB3C", X"03"),
      (X"FB3D", X"03"),
      (X"FB3E", X"03"),
      (X"FB3F", X"03"),
      (X"FB40", X"00"),
      (X"FB41", X"00"),
      (X"FB42", X"00"),
      (X"FB43", X"00"),
      (X"FB44", X"CC"),
      (X"FB45", X"CC"),
      (X"FB46", X"33"),
      (X"FB47", X"33"),
      (X"FB48", X"FF"),
      (X"FB49", X"FE"),
      (X"FB4A", X"FC"),
      (X"FB4B", X"F8"),
      (X"FB4C", X"F0"),
      (X"FB4D", X"E0"),
      (X"FB4E", X"C0"),
      (X"FB4F", X"80"),
      (X"FB50", X"03"),
      (X"FB51", X"03"),
      (X"FB52", X"03"),
      (X"FB53", X"03"),
      (X"FB54", X"03"),
      (X"FB55", X"03"),
      (X"FB56", X"03"),
      (X"FB57", X"03"),
      (X"FB58", X"18"),
      (X"FB59", X"18"),
      (X"FB5A", X"18"),
      (X"FB5B", X"1F"),
      (X"FB5C", X"1F"),
      (X"FB5D", X"18"),
      (X"FB5E", X"18"),
      (X"FB5F", X"18"),
      (X"FB60", X"00"),
      (X"FB61", X"00"),
      (X"FB62", X"00"),
      (X"FB63", X"00"),
      (X"FB64", X"0F"),
      (X"FB65", X"0F"),
      (X"FB66", X"0F"),
      (X"FB67", X"0F"),
      (X"FB68", X"18"),
      (X"FB69", X"18"),
      (X"FB6A", X"18"),
      (X"FB6B", X"1F"),
      (X"FB6C", X"1F"),
      (X"FB6D", X"00"),
      (X"FB6E", X"00"),
      (X"FB6F", X"00"),
      (X"FB70", X"00"),
      (X"FB71", X"00"),
      (X"FB72", X"00"),
      (X"FB73", X"F8"),
      (X"FB74", X"F8"),
      (X"FB75", X"18"),
      (X"FB76", X"18"),
      (X"FB77", X"18"),
      (X"FB78", X"00"),
      (X"FB79", X"00"),
      (X"FB7A", X"00"),
      (X"FB7B", X"00"),
      (X"FB7C", X"00"),
      (X"FB7D", X"00"),
      (X"FB7E", X"FF"),
      (X"FB7F", X"FF"),
      (X"FB80", X"00"),
      (X"FB81", X"00"),
      (X"FB82", X"00"),
      (X"FB83", X"1F"),
      (X"FB84", X"1F"),
      (X"FB85", X"18"),
      (X"FB86", X"18"),
      (X"FB87", X"18"),
      (X"FB88", X"18"),
      (X"FB89", X"18"),
      (X"FB8A", X"18"),
      (X"FB8B", X"FF"),
      (X"FB8C", X"FF"),
      (X"FB8D", X"00"),
      (X"FB8E", X"00"),
      (X"FB8F", X"00"),
      (X"FB90", X"00"),
      (X"FB91", X"00"),
      (X"FB92", X"00"),
      (X"FB93", X"FF"),
      (X"FB94", X"FF"),
      (X"FB95", X"18"),
      (X"FB96", X"18"),
      (X"FB97", X"18"),
      (X"FB98", X"18"),
      (X"FB99", X"18"),
      (X"FB9A", X"18"),
      (X"FB9B", X"F8"),
      (X"FB9C", X"F8"),
      (X"FB9D", X"18"),
      (X"FB9E", X"18"),
      (X"FB9F", X"18"),
      (X"FBA0", X"C0"),
      (X"FBA1", X"C0"),
      (X"FBA2", X"C0"),
      (X"FBA3", X"C0"),
      (X"FBA4", X"C0"),
      (X"FBA5", X"C0"),
      (X"FBA6", X"C0"),
      (X"FBA7", X"C0"),
      (X"FBA8", X"E0"),
      (X"FBA9", X"E0"),
      (X"FBAA", X"E0"),
      (X"FBAB", X"E0"),
      (X"FBAC", X"E0"),
      (X"FBAD", X"E0"),
      (X"FBAE", X"E0"),
      (X"FBAF", X"E0"),
      (X"FBB0", X"07"),
      (X"FBB1", X"07"),
      (X"FBB2", X"07"),
      (X"FBB3", X"07"),
      (X"FBB4", X"07"),
      (X"FBB5", X"07"),
      (X"FBB6", X"07"),
      (X"FBB7", X"07"),
      (X"FBB8", X"FF"),
      (X"FBB9", X"FF"),
      (X"FBBA", X"00"),
      (X"FBBB", X"00"),
      (X"FBBC", X"00"),
      (X"FBBD", X"00"),
      (X"FBBE", X"00"),
      (X"FBBF", X"00"),
      (X"FBC0", X"FF"),
      (X"FBC1", X"FF"),
      (X"FBC2", X"FF"),
      (X"FBC3", X"00"),
      (X"FBC4", X"00"),
      (X"FBC5", X"00"),
      (X"FBC6", X"00"),
      (X"FBC7", X"00"),
      (X"FBC8", X"00"),
      (X"FBC9", X"00"),
      (X"FBCA", X"00"),
      (X"FBCB", X"00"),
      (X"FBCC", X"00"),
      (X"FBCD", X"FF"),
      (X"FBCE", X"FF"),
      (X"FBCF", X"FF"),
      (X"FBD0", X"03"),
      (X"FBD1", X"03"),
      (X"FBD2", X"03"),
      (X"FBD3", X"03"),
      (X"FBD4", X"03"),
      (X"FBD5", X"03"),
      (X"FBD6", X"FF"),
      (X"FBD7", X"FF"),
      (X"FBD8", X"00"),
      (X"FBD9", X"00"),
      (X"FBDA", X"00"),
      (X"FBDB", X"00"),
      (X"FBDC", X"F0"),
      (X"FBDD", X"F0"),
      (X"FBDE", X"F0"),
      (X"FBDF", X"F0"),
      (X"FBE0", X"0F"),
      (X"FBE1", X"0F"),
      (X"FBE2", X"0F"),
      (X"FBE3", X"0F"),
      (X"FBE4", X"00"),
      (X"FBE5", X"00"),
      (X"FBE6", X"00"),
      (X"FBE7", X"00"),
      (X"FBE8", X"18"),
      (X"FBE9", X"18"),
      (X"FBEA", X"18"),
      (X"FBEB", X"F8"),
      (X"FBEC", X"F8"),
      (X"FBED", X"00"),
      (X"FBEE", X"00"),
      (X"FBEF", X"00"),
      (X"FBF0", X"F0"),
      (X"FBF1", X"F0"),
      (X"FBF2", X"F0"),
      (X"FBF3", X"F0"),
      (X"FBF4", X"00"),
      (X"FBF5", X"00"),
      (X"FBF6", X"00"),
      (X"FBF7", X"00"),
      (X"FBF8", X"F0"),
      (X"FBF9", X"F0"),
      (X"FBFA", X"F0"),
      (X"FBFB", X"F0"),
      (X"FBFC", X"0F"),
      (X"FBFD", X"0F"),
      (X"FBFE", X"0F"),
      (X"FBFF", X"0F"),
      (X"FC00", X"C3"),
      (X"FC01", X"99"),
      (X"FC02", X"91"),
      (X"FC03", X"91"),
      (X"FC04", X"9F"),
      (X"FC05", X"9D"),
      (X"FC06", X"C3"),
      (X"FC07", X"FF"),
      (X"FC08", X"E7"),
      (X"FC09", X"C3"),
      (X"FC0A", X"99"),
      (X"FC0B", X"81"),
      (X"FC0C", X"99"),
      (X"FC0D", X"99"),
      (X"FC0E", X"99"),
      (X"FC0F", X"FF"),
      (X"FC10", X"83"),
      (X"FC11", X"99"),
      (X"FC12", X"99"),
      (X"FC13", X"83"),
      (X"FC14", X"99"),
      (X"FC15", X"99"),
      (X"FC16", X"83"),
      (X"FC17", X"FF"),
      (X"FC18", X"C3"),
      (X"FC19", X"99"),
      (X"FC1A", X"9F"),
      (X"FC1B", X"9F"),
      (X"FC1C", X"9F"),
      (X"FC1D", X"99"),
      (X"FC1E", X"C3"),
      (X"FC1F", X"FF"),
      (X"FC20", X"87"),
      (X"FC21", X"93"),
      (X"FC22", X"99"),
      (X"FC23", X"99"),
      (X"FC24", X"99"),
      (X"FC25", X"93"),
      (X"FC26", X"87"),
      (X"FC27", X"FF"),
      (X"FC28", X"81"),
      (X"FC29", X"9F"),
      (X"FC2A", X"9F"),
      (X"FC2B", X"87"),
      (X"FC2C", X"9F"),
      (X"FC2D", X"9F"),
      (X"FC2E", X"81"),
      (X"FC2F", X"FF"),
      (X"FC30", X"81"),
      (X"FC31", X"9F"),
      (X"FC32", X"9F"),
      (X"FC33", X"87"),
      (X"FC34", X"9F"),
      (X"FC35", X"9F"),
      (X"FC36", X"9F"),
      (X"FC37", X"FF"),
      (X"FC38", X"C3"),
      (X"FC39", X"99"),
      (X"FC3A", X"9F"),
      (X"FC3B", X"91"),
      (X"FC3C", X"99"),
      (X"FC3D", X"99"),
      (X"FC3E", X"C3"),
      (X"FC3F", X"FF"),
      (X"FC40", X"99"),
      (X"FC41", X"99"),
      (X"FC42", X"99"),
      (X"FC43", X"81"),
      (X"FC44", X"99"),
      (X"FC45", X"99"),
      (X"FC46", X"99"),
      (X"FC47", X"FF"),
      (X"FC48", X"C3"),
      (X"FC49", X"E7"),
      (X"FC4A", X"E7"),
      (X"FC4B", X"E7"),
      (X"FC4C", X"E7"),
      (X"FC4D", X"E7"),
      (X"FC4E", X"C3"),
      (X"FC4F", X"FF"),
      (X"FC50", X"E1"),
      (X"FC51", X"F3"),
      (X"FC52", X"F3"),
      (X"FC53", X"F3"),
      (X"FC54", X"F3"),
      (X"FC55", X"93"),
      (X"FC56", X"C7"),
      (X"FC57", X"FF"),
      (X"FC58", X"99"),
      (X"FC59", X"93"),
      (X"FC5A", X"87"),
      (X"FC5B", X"8F"),
      (X"FC5C", X"87"),
      (X"FC5D", X"93"),
      (X"FC5E", X"99"),
      (X"FC5F", X"FF"),
      (X"FC60", X"9F"),
      (X"FC61", X"9F"),
      (X"FC62", X"9F"),
      (X"FC63", X"9F"),
      (X"FC64", X"9F"),
      (X"FC65", X"9F"),
      (X"FC66", X"81"),
      (X"FC67", X"FF"),
      (X"FC68", X"9C"),
      (X"FC69", X"88"),
      (X"FC6A", X"80"),
      (X"FC6B", X"94"),
      (X"FC6C", X"9C"),
      (X"FC6D", X"9C"),
      (X"FC6E", X"9C"),
      (X"FC6F", X"FF"),
      (X"FC70", X"99"),
      (X"FC71", X"89"),
      (X"FC72", X"81"),
      (X"FC73", X"81"),
      (X"FC74", X"91"),
      (X"FC75", X"99"),
      (X"FC76", X"99"),
      (X"FC77", X"FF"),
      (X"FC78", X"C3"),
      (X"FC79", X"99"),
      (X"FC7A", X"99"),
      (X"FC7B", X"99"),
      (X"FC7C", X"99"),
      (X"FC7D", X"99"),
      (X"FC7E", X"C3"),
      (X"FC7F", X"FF"),
      (X"FC80", X"83"),
      (X"FC81", X"99"),
      (X"FC82", X"99"),
      (X"FC83", X"83"),
      (X"FC84", X"9F"),
      (X"FC85", X"9F"),
      (X"FC86", X"9F"),
      (X"FC87", X"FF"),
      (X"FC88", X"C3"),
      (X"FC89", X"99"),
      (X"FC8A", X"99"),
      (X"FC8B", X"99"),
      (X"FC8C", X"99"),
      (X"FC8D", X"C3"),
      (X"FC8E", X"F1"),
      (X"FC8F", X"FF"),
      (X"FC90", X"83"),
      (X"FC91", X"99"),
      (X"FC92", X"99"),
      (X"FC93", X"83"),
      (X"FC94", X"87"),
      (X"FC95", X"93"),
      (X"FC96", X"99"),
      (X"FC97", X"FF"),
      (X"FC98", X"C3"),
      (X"FC99", X"99"),
      (X"FC9A", X"9F"),
      (X"FC9B", X"C3"),
      (X"FC9C", X"F9"),
      (X"FC9D", X"99"),
      (X"FC9E", X"C3"),
      (X"FC9F", X"FF"),
      (X"FCA0", X"81"),
      (X"FCA1", X"E7"),
      (X"FCA2", X"E7"),
      (X"FCA3", X"E7"),
      (X"FCA4", X"E7"),
      (X"FCA5", X"E7"),
      (X"FCA6", X"E7"),
      (X"FCA7", X"FF"),
      (X"FCA8", X"99"),
      (X"FCA9", X"99"),
      (X"FCAA", X"99"),
      (X"FCAB", X"99"),
      (X"FCAC", X"99"),
      (X"FCAD", X"99"),
      (X"FCAE", X"C3"),
      (X"FCAF", X"FF"),
      (X"FCB0", X"99"),
      (X"FCB1", X"99"),
      (X"FCB2", X"99"),
      (X"FCB3", X"99"),
      (X"FCB4", X"99"),
      (X"FCB5", X"C3"),
      (X"FCB6", X"E7"),
      (X"FCB7", X"FF"),
      (X"FCB8", X"9C"),
      (X"FCB9", X"9C"),
      (X"FCBA", X"9C"),
      (X"FCBB", X"94"),
      (X"FCBC", X"80"),
      (X"FCBD", X"88"),
      (X"FCBE", X"9C"),
      (X"FCBF", X"FF"),
      (X"FCC0", X"99"),
      (X"FCC1", X"99"),
      (X"FCC2", X"C3"),
      (X"FCC3", X"E7"),
      (X"FCC4", X"C3"),
      (X"FCC5", X"99"),
      (X"FCC6", X"99"),
      (X"FCC7", X"FF"),
      (X"FCC8", X"99"),
      (X"FCC9", X"99"),
      (X"FCCA", X"99"),
      (X"FCCB", X"C3"),
      (X"FCCC", X"E7"),
      (X"FCCD", X"E7"),
      (X"FCCE", X"E7"),
      (X"FCCF", X"FF"),
      (X"FCD0", X"81"),
      (X"FCD1", X"F9"),
      (X"FCD2", X"F3"),
      (X"FCD3", X"E7"),
      (X"FCD4", X"CF"),
      (X"FCD5", X"9F"),
      (X"FCD6", X"81"),
      (X"FCD7", X"FF"),
      (X"FCD8", X"C3"),
      (X"FCD9", X"CF"),
      (X"FCDA", X"CF"),
      (X"FCDB", X"CF"),
      (X"FCDC", X"CF"),
      (X"FCDD", X"CF"),
      (X"FCDE", X"C3"),
      (X"FCDF", X"FF"),
      (X"FCE0", X"F3"),
      (X"FCE1", X"ED"),
      (X"FCE2", X"CF"),
      (X"FCE3", X"83"),
      (X"FCE4", X"CF"),
      (X"FCE5", X"9D"),
      (X"FCE6", X"03"),
      (X"FCE7", X"FF"),
      (X"FCE8", X"C3"),
      (X"FCE9", X"F3"),
      (X"FCEA", X"F3"),
      (X"FCEB", X"F3"),
      (X"FCEC", X"F3"),
      (X"FCED", X"F3"),
      (X"FCEE", X"C3"),
      (X"FCEF", X"FF"),
      (X"FCF0", X"FF"),
      (X"FCF1", X"E7"),
      (X"FCF2", X"C3"),
      (X"FCF3", X"81"),
      (X"FCF4", X"E7"),
      (X"FCF5", X"E7"),
      (X"FCF6", X"E7"),
      (X"FCF7", X"E7"),
      (X"FCF8", X"FF"),
      (X"FCF9", X"EF"),
      (X"FCFA", X"CF"),
      (X"FCFB", X"80"),
      (X"FCFC", X"80"),
      (X"FCFD", X"CF"),
      (X"FCFE", X"EF"),
      (X"FCFF", X"FF"),
      (X"FD00", X"FF"),
      (X"FD01", X"FF"),
      (X"FD02", X"FF"),
      (X"FD03", X"FF"),
      (X"FD04", X"FF"),
      (X"FD05", X"FF"),
      (X"FD06", X"FF"),
      (X"FD07", X"FF"),
      (X"FD08", X"E7"),
      (X"FD09", X"E7"),
      (X"FD0A", X"E7"),
      (X"FD0B", X"E7"),
      (X"FD0C", X"FF"),
      (X"FD0D", X"FF"),
      (X"FD0E", X"E7"),
      (X"FD0F", X"FF"),
      (X"FD10", X"99"),
      (X"FD11", X"99"),
      (X"FD12", X"99"),
      (X"FD13", X"FF"),
      (X"FD14", X"FF"),
      (X"FD15", X"FF"),
      (X"FD16", X"FF"),
      (X"FD17", X"FF"),
      (X"FD18", X"99"),
      (X"FD19", X"99"),
      (X"FD1A", X"00"),
      (X"FD1B", X"99"),
      (X"FD1C", X"00"),
      (X"FD1D", X"99"),
      (X"FD1E", X"99"),
      (X"FD1F", X"FF"),
      (X"FD20", X"E7"),
      (X"FD21", X"C1"),
      (X"FD22", X"9F"),
      (X"FD23", X"C3"),
      (X"FD24", X"F9"),
      (X"FD25", X"83"),
      (X"FD26", X"E7"),
      (X"FD27", X"FF"),
      (X"FD28", X"9D"),
      (X"FD29", X"99"),
      (X"FD2A", X"F3"),
      (X"FD2B", X"E7"),
      (X"FD2C", X"CF"),
      (X"FD2D", X"99"),
      (X"FD2E", X"B9"),
      (X"FD2F", X"FF"),
      (X"FD30", X"C3"),
      (X"FD31", X"99"),
      (X"FD32", X"C3"),
      (X"FD33", X"C7"),
      (X"FD34", X"98"),
      (X"FD35", X"99"),
      (X"FD36", X"C0"),
      (X"FD37", X"FF"),
      (X"FD38", X"F9"),
      (X"FD39", X"F3"),
      (X"FD3A", X"E7"),
      (X"FD3B", X"FF"),
      (X"FD3C", X"FF"),
      (X"FD3D", X"FF"),
      (X"FD3E", X"FF"),
      (X"FD3F", X"FF"),
      (X"FD40", X"F3"),
      (X"FD41", X"E7"),
      (X"FD42", X"CF"),
      (X"FD43", X"CF"),
      (X"FD44", X"CF"),
      (X"FD45", X"E7"),
      (X"FD46", X"F3"),
      (X"FD47", X"FF"),
      (X"FD48", X"CF"),
      (X"FD49", X"E7"),
      (X"FD4A", X"F3"),
      (X"FD4B", X"F3"),
      (X"FD4C", X"F3"),
      (X"FD4D", X"E7"),
      (X"FD4E", X"CF"),
      (X"FD4F", X"FF"),
      (X"FD50", X"FF"),
      (X"FD51", X"99"),
      (X"FD52", X"C3"),
      (X"FD53", X"00"),
      (X"FD54", X"C3"),
      (X"FD55", X"99"),
      (X"FD56", X"FF"),
      (X"FD57", X"FF"),
      (X"FD58", X"FF"),
      (X"FD59", X"E7"),
      (X"FD5A", X"E7"),
      (X"FD5B", X"81"),
      (X"FD5C", X"E7"),
      (X"FD5D", X"E7"),
      (X"FD5E", X"FF"),
      (X"FD5F", X"FF"),
      (X"FD60", X"FF"),
      (X"FD61", X"FF"),
      (X"FD62", X"FF"),
      (X"FD63", X"FF"),
      (X"FD64", X"FF"),
      (X"FD65", X"E7"),
      (X"FD66", X"E7"),
      (X"FD67", X"CF"),
      (X"FD68", X"FF"),
      (X"FD69", X"FF"),
      (X"FD6A", X"FF"),
      (X"FD6B", X"81"),
      (X"FD6C", X"FF"),
      (X"FD6D", X"FF"),
      (X"FD6E", X"FF"),
      (X"FD6F", X"FF"),
      (X"FD70", X"FF"),
      (X"FD71", X"FF"),
      (X"FD72", X"FF"),
      (X"FD73", X"FF"),
      (X"FD74", X"FF"),
      (X"FD75", X"E7"),
      (X"FD76", X"E7"),
      (X"FD77", X"FF"),
      (X"FD78", X"FF"),
      (X"FD79", X"FC"),
      (X"FD7A", X"F9"),
      (X"FD7B", X"F3"),
      (X"FD7C", X"E7"),
      (X"FD7D", X"CF"),
      (X"FD7E", X"9F"),
      (X"FD7F", X"FF"),
      (X"FD80", X"C3"),
      (X"FD81", X"99"),
      (X"FD82", X"91"),
      (X"FD83", X"89"),
      (X"FD84", X"99"),
      (X"FD85", X"99"),
      (X"FD86", X"C3"),
      (X"FD87", X"FF"),
      (X"FD88", X"E7"),
      (X"FD89", X"E7"),
      (X"FD8A", X"C7"),
      (X"FD8B", X"E7"),
      (X"FD8C", X"E7"),
      (X"FD8D", X"E7"),
      (X"FD8E", X"81"),
      (X"FD8F", X"FF"),
      (X"FD90", X"C3"),
      (X"FD91", X"99"),
      (X"FD92", X"F9"),
      (X"FD93", X"F3"),
      (X"FD94", X"CF"),
      (X"FD95", X"9F"),
      (X"FD96", X"81"),
      (X"FD97", X"FF"),
      (X"FD98", X"C3"),
      (X"FD99", X"99"),
      (X"FD9A", X"F9"),
      (X"FD9B", X"E3"),
      (X"FD9C", X"F9"),
      (X"FD9D", X"99"),
      (X"FD9E", X"C3"),
      (X"FD9F", X"FF"),
      (X"FDA0", X"F9"),
      (X"FDA1", X"F1"),
      (X"FDA2", X"E1"),
      (X"FDA3", X"99"),
      (X"FDA4", X"80"),
      (X"FDA5", X"F9"),
      (X"FDA6", X"F9"),
      (X"FDA7", X"FF"),
      (X"FDA8", X"81"),
      (X"FDA9", X"9F"),
      (X"FDAA", X"83"),
      (X"FDAB", X"F9"),
      (X"FDAC", X"F9"),
      (X"FDAD", X"99"),
      (X"FDAE", X"C3"),
      (X"FDAF", X"FF"),
      (X"FDB0", X"C3"),
      (X"FDB1", X"99"),
      (X"FDB2", X"9F"),
      (X"FDB3", X"83"),
      (X"FDB4", X"99"),
      (X"FDB5", X"99"),
      (X"FDB6", X"C3"),
      (X"FDB7", X"FF"),
      (X"FDB8", X"81"),
      (X"FDB9", X"99"),
      (X"FDBA", X"F3"),
      (X"FDBB", X"E7"),
      (X"FDBC", X"E7"),
      (X"FDBD", X"E7"),
      (X"FDBE", X"E7"),
      (X"FDBF", X"FF"),
      (X"FDC0", X"C3"),
      (X"FDC1", X"99"),
      (X"FDC2", X"99"),
      (X"FDC3", X"C3"),
      (X"FDC4", X"99"),
      (X"FDC5", X"99"),
      (X"FDC6", X"C3"),
      (X"FDC7", X"FF"),
      (X"FDC8", X"C3"),
      (X"FDC9", X"99"),
      (X"FDCA", X"99"),
      (X"FDCB", X"C1"),
      (X"FDCC", X"F9"),
      (X"FDCD", X"99"),
      (X"FDCE", X"C3"),
      (X"FDCF", X"FF"),
      (X"FDD0", X"FF"),
      (X"FDD1", X"FF"),
      (X"FDD2", X"E7"),
      (X"FDD3", X"FF"),
      (X"FDD4", X"FF"),
      (X"FDD5", X"E7"),
      (X"FDD6", X"FF"),
      (X"FDD7", X"FF"),
      (X"FDD8", X"FF"),
      (X"FDD9", X"FF"),
      (X"FDDA", X"E7"),
      (X"FDDB", X"FF"),
      (X"FDDC", X"FF"),
      (X"FDDD", X"E7"),
      (X"FDDE", X"E7"),
      (X"FDDF", X"CF"),
      (X"FDE0", X"F1"),
      (X"FDE1", X"E7"),
      (X"FDE2", X"CF"),
      (X"FDE3", X"9F"),
      (X"FDE4", X"CF"),
      (X"FDE5", X"E7"),
      (X"FDE6", X"F1"),
      (X"FDE7", X"FF"),
      (X"FDE8", X"FF"),
      (X"FDE9", X"FF"),
      (X"FDEA", X"81"),
      (X"FDEB", X"FF"),
      (X"FDEC", X"81"),
      (X"FDED", X"FF"),
      (X"FDEE", X"FF"),
      (X"FDEF", X"FF"),
      (X"FDF0", X"8F"),
      (X"FDF1", X"E7"),
      (X"FDF2", X"F3"),
      (X"FDF3", X"F9"),
      (X"FDF4", X"F3"),
      (X"FDF5", X"E7"),
      (X"FDF6", X"8F"),
      (X"FDF7", X"FF"),
      (X"FDF8", X"C3"),
      (X"FDF9", X"99"),
      (X"FDFA", X"F9"),
      (X"FDFB", X"F3"),
      (X"FDFC", X"E7"),
      (X"FDFD", X"FF"),
      (X"FDFE", X"E7"),
      (X"FDFF", X"FF"),
      (X"FE00", X"FF"),
      (X"FE01", X"FF"),
      (X"FE02", X"FF"),
      (X"FE03", X"00"),
      (X"FE04", X"00"),
      (X"FE05", X"FF"),
      (X"FE06", X"FF"),
      (X"FE07", X"FF"),
      (X"FE08", X"F7"),
      (X"FE09", X"E3"),
      (X"FE0A", X"C1"),
      (X"FE0B", X"80"),
      (X"FE0C", X"80"),
      (X"FE0D", X"E3"),
      (X"FE0E", X"C1"),
      (X"FE0F", X"FF"),
      (X"FE10", X"E7"),
      (X"FE11", X"E7"),
      (X"FE12", X"E7"),
      (X"FE13", X"E7"),
      (X"FE14", X"E7"),
      (X"FE15", X"E7"),
      (X"FE16", X"E7"),
      (X"FE17", X"E7"),
      (X"FE18", X"FF"),
      (X"FE19", X"FF"),
      (X"FE1A", X"FF"),
      (X"FE1B", X"00"),
      (X"FE1C", X"00"),
      (X"FE1D", X"FF"),
      (X"FE1E", X"FF"),
      (X"FE1F", X"FF"),
      (X"FE20", X"FF"),
      (X"FE21", X"FF"),
      (X"FE22", X"00"),
      (X"FE23", X"00"),
      (X"FE24", X"FF"),
      (X"FE25", X"FF"),
      (X"FE26", X"FF"),
      (X"FE27", X"FF"),
      (X"FE28", X"FF"),
      (X"FE29", X"00"),
      (X"FE2A", X"00"),
      (X"FE2B", X"FF"),
      (X"FE2C", X"FF"),
      (X"FE2D", X"FF"),
      (X"FE2E", X"FF"),
      (X"FE2F", X"FF"),
      (X"FE30", X"FF"),
      (X"FE31", X"FF"),
      (X"FE32", X"FF"),
      (X"FE33", X"FF"),
      (X"FE34", X"00"),
      (X"FE35", X"00"),
      (X"FE36", X"FF"),
      (X"FE37", X"FF"),
      (X"FE38", X"CF"),
      (X"FE39", X"CF"),
      (X"FE3A", X"CF"),
      (X"FE3B", X"CF"),
      (X"FE3C", X"CF"),
      (X"FE3D", X"CF"),
      (X"FE3E", X"CF"),
      (X"FE3F", X"CF"),
      (X"FE40", X"F3"),
      (X"FE41", X"F3"),
      (X"FE42", X"F3"),
      (X"FE43", X"F3"),
      (X"FE44", X"F3"),
      (X"FE45", X"F3"),
      (X"FE46", X"F3"),
      (X"FE47", X"F3"),
      (X"FE48", X"FF"),
      (X"FE49", X"FF"),
      (X"FE4A", X"FF"),
      (X"FE4B", X"1F"),
      (X"FE4C", X"0F"),
      (X"FE4D", X"C7"),
      (X"FE4E", X"E7"),
      (X"FE4F", X"E7"),
      (X"FE50", X"E7"),
      (X"FE51", X"E7"),
      (X"FE52", X"E3"),
      (X"FE53", X"F0"),
      (X"FE54", X"F8"),
      (X"FE55", X"FF"),
      (X"FE56", X"FF"),
      (X"FE57", X"FF"),
      (X"FE58", X"E7"),
      (X"FE59", X"E7"),
      (X"FE5A", X"C7"),
      (X"FE5B", X"0F"),
      (X"FE5C", X"1F"),
      (X"FE5D", X"FF"),
      (X"FE5E", X"FF"),
      (X"FE5F", X"FF"),
      (X"FE60", X"3F"),
      (X"FE61", X"3F"),
      (X"FE62", X"3F"),
      (X"FE63", X"3F"),
      (X"FE64", X"3F"),
      (X"FE65", X"3F"),
      (X"FE66", X"00"),
      (X"FE67", X"00"),
      (X"FE68", X"3F"),
      (X"FE69", X"1F"),
      (X"FE6A", X"8F"),
      (X"FE6B", X"C7"),
      (X"FE6C", X"E3"),
      (X"FE6D", X"F1"),
      (X"FE6E", X"F8"),
      (X"FE6F", X"FC"),
      (X"FE70", X"FC"),
      (X"FE71", X"F8"),
      (X"FE72", X"F1"),
      (X"FE73", X"E3"),
      (X"FE74", X"C7"),
      (X"FE75", X"8F"),
      (X"FE76", X"1F"),
      (X"FE77", X"3F"),
      (X"FE78", X"00"),
      (X"FE79", X"00"),
      (X"FE7A", X"3F"),
      (X"FE7B", X"3F"),
      (X"FE7C", X"3F"),
      (X"FE7D", X"3F"),
      (X"FE7E", X"3F"),
      (X"FE7F", X"3F"),
      (X"FE80", X"00"),
      (X"FE81", X"00"),
      (X"FE82", X"FC"),
      (X"FE83", X"FC"),
      (X"FE84", X"FC"),
      (X"FE85", X"FC"),
      (X"FE86", X"FC"),
      (X"FE87", X"FC"),
      (X"FE88", X"FF"),
      (X"FE89", X"C3"),
      (X"FE8A", X"81"),
      (X"FE8B", X"81"),
      (X"FE8C", X"81"),
      (X"FE8D", X"81"),
      (X"FE8E", X"C3"),
      (X"FE8F", X"FF"),
      (X"FE90", X"FF"),
      (X"FE91", X"FF"),
      (X"FE92", X"FF"),
      (X"FE93", X"FF"),
      (X"FE94", X"FF"),
      (X"FE95", X"00"),
      (X"FE96", X"00"),
      (X"FE97", X"FF"),
      (X"FE98", X"C9"),
      (X"FE99", X"80"),
      (X"FE9A", X"80"),
      (X"FE9B", X"80"),
      (X"FE9C", X"C1"),
      (X"FE9D", X"E3"),
      (X"FE9E", X"F7"),
      (X"FE9F", X"FF"),
      (X"FEA0", X"9F"),
      (X"FEA1", X"9F"),
      (X"FEA2", X"9F"),
      (X"FEA3", X"9F"),
      (X"FEA4", X"9F"),
      (X"FEA5", X"9F"),
      (X"FEA6", X"9F"),
      (X"FEA7", X"9F"),
      (X"FEA8", X"FF"),
      (X"FEA9", X"FF"),
      (X"FEAA", X"FF"),
      (X"FEAB", X"F8"),
      (X"FEAC", X"F0"),
      (X"FEAD", X"E3"),
      (X"FEAE", X"E7"),
      (X"FEAF", X"E7"),
      (X"FEB0", X"3C"),
      (X"FEB1", X"18"),
      (X"FEB2", X"81"),
      (X"FEB3", X"C3"),
      (X"FEB4", X"C3"),
      (X"FEB5", X"81"),
      (X"FEB6", X"18"),
      (X"FEB7", X"3C"),
      (X"FEB8", X"FF"),
      (X"FEB9", X"C3"),
      (X"FEBA", X"81"),
      (X"FEBB", X"99"),
      (X"FEBC", X"99"),
      (X"FEBD", X"81"),
      (X"FEBE", X"C3"),
      (X"FEBF", X"FF"),
      (X"FEC0", X"E7"),
      (X"FEC1", X"E7"),
      (X"FEC2", X"99"),
      (X"FEC3", X"99"),
      (X"FEC4", X"E7"),
      (X"FEC5", X"E7"),
      (X"FEC6", X"C3"),
      (X"FEC7", X"FF"),
      (X"FEC8", X"F9"),
      (X"FEC9", X"F9"),
      (X"FECA", X"F9"),
      (X"FECB", X"F9"),
      (X"FECC", X"F9"),
      (X"FECD", X"F9"),
      (X"FECE", X"F9"),
      (X"FECF", X"F9"),
      (X"FED0", X"F7"),
      (X"FED1", X"E3"),
      (X"FED2", X"C1"),
      (X"FED3", X"80"),
      (X"FED4", X"C1"),
      (X"FED5", X"E3"),
      (X"FED6", X"F7"),
      (X"FED7", X"FF"),
      (X"FED8", X"E7"),
      (X"FED9", X"E7"),
      (X"FEDA", X"E7"),
      (X"FEDB", X"00"),
      (X"FEDC", X"00"),
      (X"FEDD", X"E7"),
      (X"FEDE", X"E7"),
      (X"FEDF", X"E7"),
      (X"FEE0", X"3F"),
      (X"FEE1", X"3F"),
      (X"FEE2", X"CF"),
      (X"FEE3", X"CF"),
      (X"FEE4", X"3F"),
      (X"FEE5", X"3F"),
      (X"FEE6", X"CF"),
      (X"FEE7", X"CF"),
      (X"FEE8", X"E7"),
      (X"FEE9", X"E7"),
      (X"FEEA", X"E7"),
      (X"FEEB", X"E7"),
      (X"FEEC", X"E7"),
      (X"FEED", X"E7"),
      (X"FEEE", X"E7"),
      (X"FEEF", X"E7"),
      (X"FEF0", X"FF"),
      (X"FEF1", X"FF"),
      (X"FEF2", X"FC"),
      (X"FEF3", X"C1"),
      (X"FEF4", X"89"),
      (X"FEF5", X"C9"),
      (X"FEF6", X"C9"),
      (X"FEF7", X"FF"),
      (X"FEF8", X"00"),
      (X"FEF9", X"80"),
      (X"FEFA", X"C0"),
      (X"FEFB", X"E0"),
      (X"FEFC", X"F0"),
      (X"FEFD", X"F8"),
      (X"FEFE", X"FC"),
      (X"FEFF", X"FE"),
      (X"FF00", X"FF"),
      (X"FF01", X"FF"),
      (X"FF02", X"FF"),
      (X"FF03", X"FF"),
      (X"FF04", X"FF"),
      (X"FF05", X"FF"),
      (X"FF06", X"FF"),
      (X"FF07", X"FF"),
      (X"FF08", X"0F"),
      (X"FF09", X"0F"),
      (X"FF0A", X"0F"),
      (X"FF0B", X"0F"),
      (X"FF0C", X"0F"),
      (X"FF0D", X"0F"),
      (X"FF0E", X"0F"),
      (X"FF0F", X"0F"),
      (X"FF10", X"FF"),
      (X"FF11", X"FF"),
      (X"FF12", X"FF"),
      (X"FF13", X"FF"),
      (X"FF14", X"00"),
      (X"FF15", X"00"),
      (X"FF16", X"00"),
      (X"FF17", X"00"),
      (X"FF18", X"00"),
      (X"FF19", X"FF"),
      (X"FF1A", X"FF"),
      (X"FF1B", X"FF"),
      (X"FF1C", X"FF"),
      (X"FF1D", X"FF"),
      (X"FF1E", X"FF"),
      (X"FF1F", X"FF"),
      (X"FF20", X"FF"),
      (X"FF21", X"FF"),
      (X"FF22", X"FF"),
      (X"FF23", X"FF"),
      (X"FF24", X"FF"),
      (X"FF25", X"FF"),
      (X"FF26", X"FF"),
      (X"FF27", X"00"),
      (X"FF28", X"3F"),
      (X"FF29", X"3F"),
      (X"FF2A", X"3F"),
      (X"FF2B", X"3F"),
      (X"FF2C", X"3F"),
      (X"FF2D", X"3F"),
      (X"FF2E", X"3F"),
      (X"FF2F", X"3F"),
      (X"FF30", X"33"),
      (X"FF31", X"33"),
      (X"FF32", X"CC"),
      (X"FF33", X"CC"),
      (X"FF34", X"33"),
      (X"FF35", X"33"),
      (X"FF36", X"CC"),
      (X"FF37", X"CC"),
      (X"FF38", X"FC"),
      (X"FF39", X"FC"),
      (X"FF3A", X"FC"),
      (X"FF3B", X"FC"),
      (X"FF3C", X"FC"),
      (X"FF3D", X"FC"),
      (X"FF3E", X"FC"),
      (X"FF3F", X"FC"),
      (X"FF40", X"FF"),
      (X"FF41", X"FF"),
      (X"FF42", X"FF"),
      (X"FF43", X"FF"),
      (X"FF44", X"33"),
      (X"FF45", X"33"),
      (X"FF46", X"CC"),
      (X"FF47", X"CC"),
      (X"FF48", X"00"),
      (X"FF49", X"01"),
      (X"FF4A", X"03"),
      (X"FF4B", X"07"),
      (X"FF4C", X"0F"),
      (X"FF4D", X"1F"),
      (X"FF4E", X"3F"),
      (X"FF4F", X"7F"),
      (X"FF50", X"FC"),
      (X"FF51", X"FC"),
      (X"FF52", X"FC"),
      (X"FF53", X"FC"),
      (X"FF54", X"FC"),
      (X"FF55", X"FC"),
      (X"FF56", X"FC"),
      (X"FF57", X"FC"),
      (X"FF58", X"E7"),
      (X"FF59", X"E7"),
      (X"FF5A", X"E7"),
      (X"FF5B", X"E0"),
      (X"FF5C", X"E0"),
      (X"FF5D", X"E7"),
      (X"FF5E", X"E7"),
      (X"FF5F", X"E7"),
      (X"FF60", X"FF"),
      (X"FF61", X"FF"),
      (X"FF62", X"FF"),
      (X"FF63", X"FF"),
      (X"FF64", X"F0"),
      (X"FF65", X"F0"),
      (X"FF66", X"F0"),
      (X"FF67", X"F0"),
      (X"FF68", X"E7"),
      (X"FF69", X"E7"),
      (X"FF6A", X"E7"),
      (X"FF6B", X"E0"),
      (X"FF6C", X"E0"),
      (X"FF6D", X"FF"),
      (X"FF6E", X"FF"),
      (X"FF6F", X"FF"),
      (X"FF70", X"FF"),
      (X"FF71", X"FF"),
      (X"FF72", X"FF"),
      (X"FF73", X"07"),
      (X"FF74", X"07"),
      (X"FF75", X"E7"),
      (X"FF76", X"E7"),
      (X"FF77", X"E7"),
      (X"FF78", X"FF"),
      (X"FF79", X"FF"),
      (X"FF7A", X"FF"),
      (X"FF7B", X"FF"),
      (X"FF7C", X"FF"),
      (X"FF7D", X"FF"),
      (X"FF7E", X"00"),
      (X"FF7F", X"00"),
      (X"FF80", X"FF"),
      (X"FF81", X"FF"),
      (X"FF82", X"FF"),
      (X"FF83", X"E0"),
      (X"FF84", X"E0"),
      (X"FF85", X"E7"),
      (X"FF86", X"E7"),
      (X"FF87", X"E7"),
      (X"FF88", X"E7"),
      (X"FF89", X"E7"),
      (X"FF8A", X"E7"),
      (X"FF8B", X"00"),
      (X"FF8C", X"00"),
      (X"FF8D", X"FF"),
      (X"FF8E", X"FF"),
      (X"FF8F", X"FF"),
      (X"FF90", X"FF"),
      (X"FF91", X"FF"),
      (X"FF92", X"FF"),
      (X"FF93", X"00"),
      (X"FF94", X"00"),
      (X"FF95", X"E7"),
      (X"FF96", X"E7"),
      (X"FF97", X"E7"),
      (X"FF98", X"E7"),
      (X"FF99", X"E7"),
      (X"FF9A", X"E7"),
      (X"FF9B", X"07"),
      (X"FF9C", X"07"),
      (X"FF9D", X"E7"),
      (X"FF9E", X"E7"),
      (X"FF9F", X"E7"),
      (X"FFA0", X"3F"),
      (X"FFA1", X"3F"),
      (X"FFA2", X"3F"),
      (X"FFA3", X"3F"),
      (X"FFA4", X"3F"),
      (X"FFA5", X"3F"),
      (X"FFA6", X"3F"),
      (X"FFA7", X"3F"),
      (X"FFA8", X"1F"),
      (X"FFA9", X"1F"),
      (X"FFAA", X"1F"),
      (X"FFAB", X"1F"),
      (X"FFAC", X"1F"),
      (X"FFAD", X"1F"),
      (X"FFAE", X"1F"),
      (X"FFAF", X"1F"),
      (X"FFB0", X"F8"),
      (X"FFB1", X"F8"),
      (X"FFB2", X"F8"),
      (X"FFB3", X"F8"),
      (X"FFB4", X"F8"),
      (X"FFB5", X"F8"),
      (X"FFB6", X"F8"),
      (X"FFB7", X"F8"),
      (X"FFB8", X"00"),
      (X"FFB9", X"00"),
      (X"FFBA", X"FF"),
      (X"FFBB", X"FF"),
      (X"FFBC", X"FF"),
      (X"FFBD", X"FF"),
      (X"FFBE", X"FF"),
      (X"FFBF", X"FF"),
      (X"FFC0", X"00"),
      (X"FFC1", X"00"),
      (X"FFC2", X"00"),
      (X"FFC3", X"FF"),
      (X"FFC4", X"FF"),
      (X"FFC5", X"FF"),
      (X"FFC6", X"FF"),
      (X"FFC7", X"FF"),
      (X"FFC8", X"FF"),
      (X"FFC9", X"FF"),
      (X"FFCA", X"FF"),
      (X"FFCB", X"FF"),
      (X"FFCC", X"FF"),
      (X"FFCD", X"00"),
      (X"FFCE", X"00"),
      (X"FFCF", X"00"),
      (X"FFD0", X"FC"),
      (X"FFD1", X"FC"),
      (X"FFD2", X"FC"),
      (X"FFD3", X"FC"),
      (X"FFD4", X"FC"),
      (X"FFD5", X"FC"),
      (X"FFD6", X"00"),
      (X"FFD7", X"00"),
      (X"FFD8", X"FF"),
      (X"FFD9", X"FF"),
      (X"FFDA", X"FF"),
      (X"FFDB", X"FF"),
      (X"FFDC", X"0F"),
      (X"FFDD", X"0F"),
      (X"FFDE", X"0F"),
      (X"FFDF", X"0F"),
      (X"FFE0", X"F0"),
      (X"FFE1", X"F0"),
      (X"FFE2", X"F0"),
      (X"FFE3", X"F0"),
      (X"FFE4", X"FF"),
      (X"FFE5", X"FF"),
      (X"FFE6", X"FF"),
      (X"FFE7", X"FF"),
      (X"FFE8", X"E7"),
      (X"FFE9", X"E7"),
      (X"FFEA", X"E7"),
      (X"FFEB", X"07"),
      (X"FFEC", X"07"),
      (X"FFED", X"FF"),
      (X"FFEE", X"FF"),
      (X"FFEF", X"FF"),
      (X"FFF0", X"0F"),
      (X"FFF1", X"0F"),
      (X"FFF2", X"0F"),
      (X"FFF3", X"0F"),
      (X"FFF4", X"FF"),
      (X"FFF5", X"FF"),
      (X"FFF6", X"FF"),
      (X"FFF7", X"FF"),
      (X"FFF8", X"0F"),
      (X"FFF9", X"0F"),
      (X"FFFA", X"0F"),
      (X"FFFB", X"0F"),
      (X"FFFC", X"F0"),
      (X"FFFD", X"F0"),
      (X"FFFE", X"F0"),
      (X"FFFF", X"F0")
   );

   signal wr_index : integer := 0;

begin

   -- This is a temporary process that populates the VRAM
   p_wr : process (clk_i)
   begin
      if rising_edge(clk_i) then
         wr_en_o <= '0';
         if wr_index < wr_default'length then
            wr_addr_o <= "0" & wr_default(wr_index).addr;
            wr_en_o   <= '1';
            wr_data_o <= wr_default(wr_index).data;
            wr_index  <= wr_index + 1;
         end if;
      end if;
   end process p_wr;

end architecture structural;


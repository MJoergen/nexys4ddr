--------------------------------------
-- The Control Logic
--

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ctl is
   port (
      clk_i  : in  std_logic;
      rst_i  : in  std_logic;
      data_i : in  std_logic_vector( 7 downto 0);

      mem_rden_o      : out std_logic;    -- Read from memory
      mem_wren_o      : out std_logic;    -- Write to memory
      mem_addr_wren_o : out std_logic;    -- Write to address hold register
      mem_addr_sel_o  : out std_logic_vector(1 downto 0);   -- Memory address select
      mem_data_sel_o  : out std_logic_vector(1 downto 0);   -- Memory data select
      reg_wren_o      : out std_logic;    -- Write to register file
      reg_nr_o        : out std_logic_vector(1 downto 0);   -- Register number
      pc_sel_o        : out std_logic_vector(1 downto 0);   -- PC relect
      alu_func_o      : out std_logic_vector(3 downto 0);   -- ALU function
      clc_o           : out std_logic;                      -- Clear carry
      sr_alu_wren_o   : out std_logic;                      -- Write status register
      sp_sel_o        : out std_logic_vector(1 downto 0);   -- Stack pointer update

      debug_o : out std_logic_vector(10 downto 0)
   );
end ctl;

architecture Structural of ctl is

   signal cnt_r   : std_logic_vector(2 downto 0) := (others => '0');
   signal inst_r  : std_logic_vector(7 downto 0) := (others => '0');
   signal last    : std_logic;
   signal invalid : std_logic;

   signal ctl     : std_logic_vector(21 downto 0);

begin

   mem_rden_o      <= ctl(0);
   mem_wren_o      <= ctl(1);
   mem_addr_wren_o <= ctl(2);
   mem_addr_sel_o  <= ctl(4 downto 3);
   mem_data_sel_o  <= ctl(6 downto 5);
   reg_wren_o      <= ctl(7);
   reg_nr_o        <= ctl(9 downto 8);
   pc_sel_o        <= ctl(11 downto 10);
   alu_func_o      <= ctl(15 downto 12);
   clc_o           <= ctl(16);
   sr_alu_wren_o   <= ctl(17);
   last            <= ctl(18);
   invalid         <= ctl(19);
   sp_sel_o        <= ctl(21 downto 20);

   p_assert : process (clk_i)
   begin 
      if rising_edge(clk_i) then
         assert rst_i /= '0' or invalid = '0' report "Invalid opcode" severity failure;
      end if;
   end process p_assert;

   debug_o( 7 downto 0) <= inst_r;
   debug_o(10 downto 8) <= cnt_r;

   -- Store the microinstruction counter
   p_cnt : process (clk_i)
   begin
      if rising_edge(clk_i) then
         cnt_r <= cnt_r + 1;

         if rst_i = '1' or last = '1' then
            cnt_r <= (others => '0');
         end if;
      end if;
   end process p_cnt;


   -- Store the current instruction
   p_inst : process (clk_i)
   begin
      if rising_edge(clk_i) then
         if cnt_r = 0 then
            inst_r <= data_i;
         end if;
      end if;
   end process p_inst;


   -- Combinatorial process
   process (cnt_r, inst_r)
   begin
      ctl <= "0000000000000000000000";  -- Default value to avoid latch.

      if cnt_r = 0 then
         ctl <= "0000000000000000000001";
      end if;

      if cnt_r = 1 then
         case inst_r is
            when "00000000" => ctl <= B"10_0_0_0_0_0000_00_00_0_01_10_0_1_0";
            when "00000001" => ctl <= B"00_1000000000000000000_0";
            when "00000010" => ctl <= B"00_1000000000000000000_0";
            when "00000011" => ctl <= B"00_1000000000000000000_0";
            when "00000100" => ctl <= B"00_1000000000000000000_0";
            when "00000101" => ctl <= B"00_0000000000000000010_1";
            when "00000110" => ctl <= B"00_1000000000000000000_0";
            when "00000111" => ctl <= B"00_1000000000000000000_0";
            when "00001000" => ctl <= B"00_1000000000000000000_0";
            when "00001001" => ctl <= B"00_0110000000001000000_1"; -- 09 ORA #
            when "00001010" => ctl <= B"00_1000000000000000000_0";
            when "00001011" => ctl <= B"00_1000000000000000000_0";
            when "00001100" => ctl <= B"00_1000000000000000000_0";
            when "00001101" => ctl <= B"00_1000000000000000000_0";
            when "00001110" => ctl <= B"00_1000000000000000000_0";
            when "00001111" => ctl <= B"00_1000000000000000000_0";

            when "00010000" => ctl <= B"00_1000000000000000000_0";
            when "00010001" => ctl <= B"00_1000000000000000000_0";
            when "00010010" => ctl <= B"00_1000000000000000000_0";
            when "00010011" => ctl <= B"00_1000000000000000000_0";
            when "00010100" => ctl <= B"00_1000000000000000000_0";
            when "00010101" => ctl <= B"00_0000000000000000010_1";
            when "00010110" => ctl <= B"00_1000000000000000000_0";
            when "00010111" => ctl <= B"00_1000000000000000000_0";
            when "00011000" => ctl <= B"00_0101000011000000000_0";
            when "00011001" => ctl <= B"00_1000000000000000000_0";
            when "00011010" => ctl <= B"00_1000000000000000000_0";
            when "00011011" => ctl <= B"00_1000000000000000000_0";
            when "00011100" => ctl <= B"00_1000000000000000000_0";
            when "00011101" => ctl <= B"00_1000000000000000000_0";
            when "00011110" => ctl <= B"00_1000000000000000000_0";
            when "00011111" => ctl <= B"00_1000000000000000000_0";

            when "00100000" => ctl <= B"00_1000000000000000000_0";
            when "00100001" => ctl <= B"00_1000000000000000000_0";
            when "00100010" => ctl <= B"00_1000000000000000000_0";
            when "00100011" => ctl <= B"00_1000000000000000000_0";
            when "00100100" => ctl <= B"00_1000000000000000000_0";
            when "00100101" => ctl <= B"00_1000000000000000000_0";
            when "00100110" => ctl <= B"00_1000000000000000000_0";
            when "00100111" => ctl <= B"00_1000000000000000000_0";
            when "00101000" => ctl <= B"00_1000000000000000000_0";
            when "00101001" => ctl <= B"00_0110000100001000000_1"; -- 29 AND #
            when "00101010" => ctl <= B"00_1000000000000000000_0";
            when "00101011" => ctl <= B"00_1000000000000000000_0";
            when "00101100" => ctl <= B"00_1000000000000000000_0";
            when "00101101" => ctl <= B"00_1000000000000000000_0";
            when "00101110" => ctl <= B"00_1000000000000000000_0";
            when "00101111" => ctl <= B"00_1000000000000000000_0";

            when "00110000" => ctl <= B"00_1000000000000000000_0";
            when "00110001" => ctl <= B"00_1000000000000000000_0";
            when "00110010" => ctl <= B"00_1000000000000000000_0";
            when "00110011" => ctl <= B"00_1000000000000000000_0";
            when "00110100" => ctl <= B"00_1000000000000000000_0";
            when "00110101" => ctl <= B"00_1000000000000000000_0";
            when "00110110" => ctl <= B"00_1000000000000000000_0";
            when "00110111" => ctl <= B"00_1000000000000000000_0";
            when "00111000" => ctl <= B"00_1000000000000000000_0";
            when "00111001" => ctl <= B"00_1000000000000000000_0";
            when "00111010" => ctl <= B"00_1000000000000000000_0";
            when "00111011" => ctl <= B"00_1000000000000000000_0";
            when "00111100" => ctl <= B"00_1000000000000000000_0";
            when "00111101" => ctl <= B"00_1000000000000000000_0";
            when "00111110" => ctl <= B"00_1000000000000000000_0";
            when "00111111" => ctl <= B"00_1000000000000000000_0";

            when "01000000" => ctl <= B"00_1000000000000000000_0";
            when "01000001" => ctl <= B"00_1000000000000000000_0";
            when "01000010" => ctl <= B"00_1000000000000000000_0";
            when "01000011" => ctl <= B"00_1000000000000000000_0";
            when "01000100" => ctl <= B"00_1000000000000000000_0";
            when "01000101" => ctl <= B"00_0000000000000000010_1";
            when "01000110" => ctl <= B"00_1000000000000000000_0";
            when "01000111" => ctl <= B"00_1000000000000000000_0";
            when "01001000" => ctl <= B"00_1000000000000000000_0";
            when "01001001" => ctl <= B"00_0110001000001000000_1"; -- 49 EOR #
            when "01001010" => ctl <= B"00_1000000000000000000_0";
            when "01001011" => ctl <= B"00_1000000000000000000_0";
            when "01001100" => ctl <= B"00_0000000000000000010_1";
            when "01001101" => ctl <= B"00_1000000000000000000_0";
            when "01001110" => ctl <= B"00_1000000000000000000_0";
            when "01001111" => ctl <= B"00_1000000000000000000_0";

            when "01010000" => ctl <= B"00_1000000000000000000_0";
            when "01010001" => ctl <= B"00_1000000000000000000_0";
            when "01010010" => ctl <= B"00_1000000000000000000_0";
            when "01010011" => ctl <= B"00_1000000000000000000_0";
            when "01010100" => ctl <= B"00_1000000000000000000_0";
            when "01010101" => ctl <= B"00_1000000000000000000_0";
            when "01010110" => ctl <= B"00_1000000000000000000_0";
            when "01010111" => ctl <= B"00_1000000000000000000_0";
            when "01011000" => ctl <= B"00_1000000000000000000_0";
            when "01011001" => ctl <= B"00_1000000000000000000_0";
            when "01011010" => ctl <= B"00_1000000000000000000_0";
            when "01011011" => ctl <= B"00_1000000000000000000_0";
            when "01011100" => ctl <= B"00_1000000000000000000_0";
            when "01011101" => ctl <= B"00_1000000000000000000_0";
            when "01011110" => ctl <= B"00_1000000000000000000_0";
            when "01011111" => ctl <= B"00_1000000000000000000_0";

            when "01100000" => ctl <= B"00_1000000000000000000_0";
            when "01100001" => ctl <= B"00_1000000000000000000_0";
            when "01100010" => ctl <= B"00_1000000000000000000_0";
            when "01100011" => ctl <= B"00_1000000000000000000_0";
            when "01100100" => ctl <= B"00_1000000000000000000_0";
            when "01100101" => ctl <= B"00_0000000000000000010_1";
            when "01100110" => ctl <= B"00_1000000000000000000_0";
            when "01100111" => ctl <= B"00_1000000000000000000_0";
            when "01101000" => ctl <= B"00_1000000000000000000_0";
            when "01101001" => ctl <= B"00_0110001100001000000_1"; -- 69 ADC #
            when "01101010" => ctl <= B"00_1000000000000000000_0";
            when "01101011" => ctl <= B"00_1000000000000000000_0";
            when "01101100" => ctl <= B"00_1000000000000000000_0";
            when "01101101" => ctl <= B"00_1000000000000000000_0";
            when "01101110" => ctl <= B"00_1000000000000000000_0";
            when "01101111" => ctl <= B"00_1000000000000000000_0";

            when "01110000" => ctl <= B"00_1000000000000000000_0";
            when "01110001" => ctl <= B"00_1000000000000000000_0";
            when "01110010" => ctl <= B"00_1000000000000000000_0";
            when "01110011" => ctl <= B"00_1000000000000000000_0";
            when "01110100" => ctl <= B"00_1000000000000000000_0";
            when "01110101" => ctl <= B"00_1000000000000000000_0";
            when "01110110" => ctl <= B"00_1000000000000000000_0";
            when "01110111" => ctl <= B"00_1000000000000000000_0";
            when "01111000" => ctl <= B"00_1000000000000000000_0";
            when "01111001" => ctl <= B"00_1000000000000000000_0";
            when "01111010" => ctl <= B"00_1000000000000000000_0";
            when "01111011" => ctl <= B"00_1000000000000000000_0";
            when "01111100" => ctl <= B"00_1000000000000000000_0";
            when "01111101" => ctl <= B"00_1000000000000000000_0";
            when "01111110" => ctl <= B"00_1000000000000000000_0";
            when "01111111" => ctl <= B"00_1000000000000000000_0";

            when "10000000" => ctl <= B"00_1000000000000000000_0";
            when "10000001" => ctl <= B"00_1000000000000000000_0";
            when "10000010" => ctl <= B"00_1000000000000000000_0";
            when "10000011" => ctl <= B"00_1000000000000000000_0";
            when "10000100" => ctl <= B"00_1000000000000000000_0";
            when "10000101" => ctl <= B"00_0000000000000000010_1";
            when "10000110" => ctl <= B"00_1000000000000000000_0";
            when "10000111" => ctl <= B"00_1000000000000000000_0";
            when "10001000" => ctl <= B"00_1000000000000000000_0";
            when "10001001" => ctl <= B"00_1000000000000000000_0";
            when "10001010" => ctl <= B"00_1000000000000000000_0";
            when "10001011" => ctl <= B"00_1000000000000000000_0";
            when "10001100" => ctl <= B"00_1000000000000000000_0";
            when "10001101" => ctl <= B"00_1000000000000000000_0";
            when "10001110" => ctl <= B"00_1000000000000000000_0";
            when "10001111" => ctl <= B"00_1000000000000000000_0";

            when "10010000" => ctl <= B"00_1000000000000000000_0";
            when "10010001" => ctl <= B"00_1000000000000000000_0";
            when "10010010" => ctl <= B"00_1000000000000000000_0";
            when "10010011" => ctl <= B"00_1000000000000000000_0";
            when "10010100" => ctl <= B"00_1000000000000000000_0";
            when "10010101" => ctl <= B"00_1000000000000000000_0";
            when "10010110" => ctl <= B"00_1000000000000000000_0";
            when "10010111" => ctl <= B"00_1000000000000000000_0";
            when "10011000" => ctl <= B"00_1000000000000000000_0";
            when "10011001" => ctl <= B"00_1000000000000000000_0";
            when "10011010" => ctl <= B"00_1000000000000000000_0";
            when "10011011" => ctl <= B"00_1000000000000000000_0";
            when "10011100" => ctl <= B"00_1000000000000000000_0";
            when "10011101" => ctl <= B"00_1000000000000000000_0";
            when "10011110" => ctl <= B"00_1000000000000000000_0";
            when "10011111" => ctl <= B"00_1000000000000000000_0";

            when "10100000" => ctl <= B"00_1000000000000000000_0";
            when "10100001" => ctl <= B"00_1000000000000000000_0";
            when "10100010" => ctl <= B"00_1000000000000000000_0";
            when "10100011" => ctl <= B"00_1000000000000000000_0";
            when "10100100" => ctl <= B"00_1000000000000000000_0";
            when "10100101" => ctl <= B"00_0000000000000000010_1";
            when "10100110" => ctl <= B"00_1000000000000000000_0";
            when "10100111" => ctl <= B"00_1000000000000000000_0";
            when "10101000" => ctl <= B"00_1000000000000000000_0";
            when "10101001" => ctl <= B"00_0110010100001000000_1"; -- A9 LDA #
            when "10101010" => ctl <= B"00_1000000000000000000_0";
            when "10101011" => ctl <= B"00_1000000000000000000_0";
            when "10101100" => ctl <= B"00_1000000000000000000_0";
            when "10101101" => ctl <= B"00_1000000000000000000_0";
            when "10101110" => ctl <= B"00_1000000000000000000_0";
            when "10101111" => ctl <= B"00_1000000000000000000_0";

            when "10110000" => ctl <= B"00_1000000000000000000_0";
            when "10110001" => ctl <= B"00_1000000000000000000_0";
            when "10110010" => ctl <= B"00_1000000000000000000_0";
            when "10110011" => ctl <= B"00_1000000000000000000_0";
            when "10110100" => ctl <= B"00_1000000000000000000_0";
            when "10110101" => ctl <= B"00_1000000000000000000_0";
            when "10110110" => ctl <= B"00_1000000000000000000_0";
            when "10110111" => ctl <= B"00_1000000000000000000_0";
            when "10111000" => ctl <= B"00_1000000000000000000_0";
            when "10111001" => ctl <= B"00_1000000000000000000_0";
            when "10111010" => ctl <= B"00_1000000000000000000_0";
            when "10111011" => ctl <= B"00_1000000000000000000_0";
            when "10111100" => ctl <= B"00_1000000000000000000_0";
            when "10111101" => ctl <= B"00_1000000000000000000_0";
            when "10111110" => ctl <= B"00_1000000000000000000_0";
            when "10111111" => ctl <= B"00_1000000000000000000_0";

            when "11000000" => ctl <= B"00_1000000000000000000_0";
            when "11000001" => ctl <= B"00_1000000000000000000_0";
            when "11000010" => ctl <= B"00_1000000000000000000_0";
            when "11000011" => ctl <= B"00_1000000000000000000_0";
            when "11000100" => ctl <= B"00_1000000000000000000_0";
            when "11000101" => ctl <= B"00_0000000000000000010_1";
            when "11000110" => ctl <= B"00_1000000000000000000_0";
            when "11000111" => ctl <= B"00_1000000000000000000_0";
            when "11001000" => ctl <= B"00_1000000000000000000_0";
            when "11001001" => ctl <= B"00_0110011000001000000_1"; -- C9 CMP #
            when "11001010" => ctl <= B"00_1000000000000000000_0";
            when "11001011" => ctl <= B"00_1000000000000000000_0";
            when "11001100" => ctl <= B"00_1000000000000000000_0";
            when "11001101" => ctl <= B"00_1000000000000000000_0";
            when "11001110" => ctl <= B"00_1000000000000000000_0";
            when "11001111" => ctl <= B"00_1000000000000000000_0";

            when "11010000" => ctl <= B"00_1000000000000000000_0";
            when "11010001" => ctl <= B"00_1000000000000000000_0";
            when "11010010" => ctl <= B"00_1000000000000000000_0";
            when "11010011" => ctl <= B"00_1000000000000000000_0";
            when "11010100" => ctl <= B"00_1000000000000000000_0";
            when "11010101" => ctl <= B"00_1000000000000000000_0";
            when "11010110" => ctl <= B"00_1000000000000000000_0";
            when "11010111" => ctl <= B"00_1000000000000000000_0";
            when "11011000" => ctl <= B"00_1000000000000000000_0";
            when "11011001" => ctl <= B"00_1000000000000000000_0";
            when "11011010" => ctl <= B"00_1000000000000000000_0";
            when "11011011" => ctl <= B"00_1000000000000000000_0";
            when "11011100" => ctl <= B"00_1000000000000000000_0";
            when "11011101" => ctl <= B"00_1000000000000000000_0";
            when "11011110" => ctl <= B"00_1000000000000000000_0";
            when "11011111" => ctl <= B"00_1000000000000000000_0";

            when "11100000" => ctl <= B"00_1000000000000000000_0";
            when "11100001" => ctl <= B"00_1000000000000000000_0";
            when "11100010" => ctl <= B"00_1000000000000000000_0";
            when "11100011" => ctl <= B"00_1000000000000000000_0";
            when "11100100" => ctl <= B"00_1000000000000000000_0";
            when "11100101" => ctl <= B"00_0000000000000000010_1";
            when "11100110" => ctl <= B"00_1000000000000000000_0";
            when "11100111" => ctl <= B"00_1000000000000000000_0";
            when "11101000" => ctl <= B"00_1000000000000000000_0";
            when "11101001" => ctl <= B"00_0110011100001000000_1"; -- E9 SBC #
            when "11101010" => ctl <= B"00_1000000000000000000_0";
            when "11101011" => ctl <= B"00_1000000000000000000_0";
            when "11101100" => ctl <= B"00_1000000000000000000_0";
            when "11101101" => ctl <= B"00_1000000000000000000_0";
            when "11101110" => ctl <= B"00_1000000000000000000_0";
            when "11101111" => ctl <= B"00_1000000000000000000_0";

            when "11110000" => ctl <= B"00_1000000000000000000_0";
            when "11110001" => ctl <= B"00_1000000000000000000_0";
            when "11110010" => ctl <= B"00_1000000000000000000_0";
            when "11110011" => ctl <= B"00_1000000000000000000_0";
            when "11110100" => ctl <= B"00_1000000000000000000_0";
            when "11110101" => ctl <= B"00_1000000000000000000_0";
            when "11110110" => ctl <= B"00_1000000000000000000_0";
            when "11110111" => ctl <= B"00_1000000000000000000_0";
            when "11111000" => ctl <= B"00_1000000000000000000_0";
            when "11111001" => ctl <= B"00_1000000000000000000_0";
            when "11111010" => ctl <= B"00_1000000000000000000_0";
            when "11111011" => ctl <= B"00_1000000000000000000_0";
            when "11111100" => ctl <= B"00_1000000000000000000_0";
            when "11111101" => ctl <= B"00_1000000000000000000_0";
            when "11111110" => ctl <= B"00_1000000000000000000_0";
            when "11111111" => ctl <= B"00_1000000000000000000_0";

            -- Default to avoid latch
            when others => ctl <= "0010000000000000000000";
         end case;
      end if;

      if cnt_r = 2 then
         case inst_r is
            when "00000000" => ctl <= "1000000000000001010010";
            when "00000001" => ctl <= "0010000000000000000000";
            when "00000010" => ctl <= "0010000000000000000000";
            when "00000011" => ctl <= "0010000000000000000000";
            when "00000100" => ctl <= "0010000000000000000000";
            when "00000101" => ctl <= "0001100000110010001001";
            when "00000110" => ctl <= "0010000000000000000000";
            when "00000111" => ctl <= "0010000000000000000000";
            when "00001000" => ctl <= "0010000000000000000000";
            when "00001001" => ctl <= "0010000000000000000000";
            when "00001010" => ctl <= "0010000000000000000000";
            when "00001011" => ctl <= "0010000000000000000000";
            when "00001100" => ctl <= "0010000000000000000000";
            when "00001101" => ctl <= "0010000000000000000000";
            when "00001110" => ctl <= "0010000000000000000000";
            when "00001111" => ctl <= "0010000000000000000000";

            when "00010000" => ctl <= "0010000000000000000000";
            when "00010001" => ctl <= "0010000000000000000000";
            when "00010010" => ctl <= "0010000000000000000000";
            when "00010011" => ctl <= "0010000000000000000000";
            when "00010100" => ctl <= "0010000000000000000000";
            when "00010101" => ctl <= "0010000000000000000000";
            when "00010110" => ctl <= "0010000000000000000000";
            when "00010111" => ctl <= "0010000000000000000000";
            when "00011000" => ctl <= "0010000000000000000000";
            when "00011001" => ctl <= "0010000000000000000000";
            when "00011010" => ctl <= "0010000000000000000000";
            when "00011011" => ctl <= "0010000000000000000000";
            when "00011100" => ctl <= "0010000000000000000000";
            when "00011101" => ctl <= "0010000000000000000000";
            when "00011110" => ctl <= "0010000000000000000000";
            when "00011111" => ctl <= "0010000000000000000000";

            when "00100000" => ctl <= "0010000000000000000000";
            when "00100001" => ctl <= "0010000000000000000000";
            when "00100010" => ctl <= "0010000000000000000000";
            when "00100011" => ctl <= "0010000000000000000000";
            when "00100100" => ctl <= "0010000000000000000000";
            when "00100101" => ctl <= "0001100001110010001001";
            when "00100110" => ctl <= "0010000000000000000000";
            when "00100111" => ctl <= "0010000000000000000000";
            when "00101000" => ctl <= "0010000000000000000000";
            when "00101001" => ctl <= "0010000000000000000000";
            when "00101010" => ctl <= "0010000000000000000000";
            when "00101011" => ctl <= "0010000000000000000000";
            when "00101100" => ctl <= "0010000000000000000000";
            when "00101101" => ctl <= "0010000000000000000000";
            when "00101110" => ctl <= "0010000000000000000000";
            when "00101111" => ctl <= "0010000000000000000000";

            when "00110000" => ctl <= "0010000000000000000000";
            when "00110001" => ctl <= "0010000000000000000000";
            when "00110010" => ctl <= "0010000000000000000000";
            when "00110011" => ctl <= "0010000000000000000000";
            when "00110100" => ctl <= "0010000000000000000000";
            when "00110101" => ctl <= "0010000000000000000000";
            when "00110110" => ctl <= "0010000000000000000000";
            when "00110111" => ctl <= "0010000000000000000000";
            when "00111000" => ctl <= "0010000000000000000000";
            when "00111001" => ctl <= "0010000000000000000000";
            when "00111010" => ctl <= "0010000000000000000000";
            when "00111011" => ctl <= "0010000000000000000000";
            when "00111100" => ctl <= "0010000000000000000000";
            when "00111101" => ctl <= "0010000000000000000000";
            when "00111110" => ctl <= "0010000000000000000000";
            when "00111111" => ctl <= "0010000000000000000000";

            when "01000000" => ctl <= "0010000000000000000000";
            when "01000001" => ctl <= "0010000000000000000000";
            when "01000010" => ctl <= "0010000000000000000000";
            when "01000011" => ctl <= "0010000000000000000000";
            when "01000100" => ctl <= "0010000000000000000000";
            when "01000101" => ctl <= "0001100010110010001001";
            when "01000110" => ctl <= "0010000000000000000000";
            when "01000111" => ctl <= "0010000000000000000000";
            when "01001000" => ctl <= "0010000000000000000000";
            when "01001001" => ctl <= "0010000000000000000000";
            when "01001010" => ctl <= "0010000000000000000000";
            when "01001011" => ctl <= "0010000000000000000000";
            when "01001100" => ctl <= "0001000000010000000001";
            when "01001101" => ctl <= "0010000000000000000000";
            when "01001110" => ctl <= "0010000000000000000000";
            when "01001111" => ctl <= "0010000000000000000000";

            when "01010000" => ctl <= "0010000000000000000000";
            when "01010001" => ctl <= "0010000000000000000000";
            when "01010010" => ctl <= "0010000000000000000000";
            when "01010011" => ctl <= "0010000000000000000000";
            when "01010100" => ctl <= "0010000000000000000000";
            when "01010101" => ctl <= "0010000000000000000000";
            when "01010110" => ctl <= "0010000000000000000000";
            when "01010111" => ctl <= "0010000000000000000000";
            when "01011000" => ctl <= "0010000000000000000000";
            when "01011001" => ctl <= "0010000000000000000000";
            when "01011010" => ctl <= "0010000000000000000000";
            when "01011011" => ctl <= "0010000000000000000000";
            when "01011100" => ctl <= "0010000000000000000000";
            when "01011101" => ctl <= "0010000000000000000000";
            when "01011110" => ctl <= "0010000000000000000000";
            when "01011111" => ctl <= "0010000000000000000000";

            when "01100000" => ctl <= "0010000000000000000000";
            when "01100001" => ctl <= "0010000000000000000000";
            when "01100010" => ctl <= "0010000000000000000000";
            when "01100011" => ctl <= "0010000000000000000000";
            when "01100100" => ctl <= "0010000000000000000000";
            when "01100101" => ctl <= "0001100011110010001001";
            when "01100110" => ctl <= "0010000000000000000000";
            when "01100111" => ctl <= "0010000000000000000000";
            when "01101000" => ctl <= "0010000000000000000000";
            when "01101001" => ctl <= "0010000000000000000000";
            when "01101010" => ctl <= "0010000000000000000000";
            when "01101011" => ctl <= "0010000000000000000000";
            when "01101100" => ctl <= "0010000000000000000000";
            when "01101101" => ctl <= "0010000000000000000000";
            when "01101110" => ctl <= "0010000000000000000000";
            when "01101111" => ctl <= "0010000000000000000000";

            when "01110000" => ctl <= "0010000000000000000000";
            when "01110001" => ctl <= "0010000000000000000000";
            when "01110010" => ctl <= "0010000000000000000000";
            when "01110011" => ctl <= "0010000000000000000000";
            when "01110100" => ctl <= "0010000000000000000000";
            when "01110101" => ctl <= "0010000000000000000000";
            when "01110110" => ctl <= "0010000000000000000000";
            when "01110111" => ctl <= "0010000000000000000000";
            when "01111000" => ctl <= "0010000000000000000000";
            when "01111001" => ctl <= "0010000000000000000000";
            when "01111010" => ctl <= "0010000000000000000000";
            when "01111011" => ctl <= "0010000000000000000000";
            when "01111100" => ctl <= "0010000000000000000000";
            when "01111101" => ctl <= "0010000000000000000000";
            when "01111110" => ctl <= "0010000000000000000000";
            when "01111111" => ctl <= "0010000000000000000000";

            when "10000000" => ctl <= "0010000000000000000000";
            when "10000001" => ctl <= "0010000000000000000000";
            when "10000010" => ctl <= "0010000000000000000000";
            when "10000011" => ctl <= "0010000000000000000000";
            when "10000100" => ctl <= "0010000000000000000000";
            when "10000101" => ctl <= "0001100100110010001010";
            when "10000110" => ctl <= "0010000000000000000000";
            when "10000111" => ctl <= "0010000000000000000000";
            when "10001000" => ctl <= "0010000000000000000000";
            when "10001001" => ctl <= "0010000000000000000000";
            when "10001010" => ctl <= "0010000000000000000000";
            when "10001011" => ctl <= "0010000000000000000000";
            when "10001100" => ctl <= "0010000000000000000000";
            when "10001101" => ctl <= "0010000000000000000000";
            when "10001110" => ctl <= "0010000000000000000000";
            when "10001111" => ctl <= "0010000000000000000000";

            when "10010000" => ctl <= "0010000000000000000000";
            when "10010001" => ctl <= "0010000000000000000000";
            when "10010010" => ctl <= "0010000000000000000000";
            when "10010011" => ctl <= "0010000000000000000000";
            when "10010100" => ctl <= "0010000000000000000000";
            when "10010101" => ctl <= "0010000000000000000000";
            when "10010110" => ctl <= "0010000000000000000000";
            when "10010111" => ctl <= "0010000000000000000000";
            when "10011000" => ctl <= "0010000000000000000000";
            when "10011001" => ctl <= "0010000000000000000000";
            when "10011010" => ctl <= "0010000000000000000000";
            when "10011011" => ctl <= "0010000000000000000000";
            when "10011100" => ctl <= "0010000000000000000000";
            when "10011101" => ctl <= "0010000000000000000000";
            when "10011110" => ctl <= "0010000000000000000000";
            when "10011111" => ctl <= "0010000000000000000000";

            when "10100000" => ctl <= "0010000000000000000000";
            when "10100001" => ctl <= "0010000000000000000000";
            when "10100010" => ctl <= "0010000000000000000000";
            when "10100011" => ctl <= "0010000000000000000000";
            when "10100100" => ctl <= "0010000000000000000000";
            when "10100101" => ctl <= "0001100101110010001001";
            when "10100110" => ctl <= "0010000000000000000000";
            when "10100111" => ctl <= "0010000000000000000000";
            when "10101000" => ctl <= "0010000000000000000000";
            when "10101001" => ctl <= "0010000000000000000000";
            when "10101010" => ctl <= "0010000000000000000000";
            when "10101011" => ctl <= "0010000000000000000000";
            when "10101100" => ctl <= "0010000000000000000000";
            when "10101101" => ctl <= "0010000000000000000000";
            when "10101110" => ctl <= "0010000000000000000000";
            when "10101111" => ctl <= "0010000000000000000000";

            when "10110000" => ctl <= "0010000000000000000000";
            when "10110001" => ctl <= "0010000000000000000000";
            when "10110010" => ctl <= "0010000000000000000000";
            when "10110011" => ctl <= "0010000000000000000000";
            when "10110100" => ctl <= "0010000000000000000000";
            when "10110101" => ctl <= "0010000000000000000000";
            when "10110110" => ctl <= "0010000000000000000000";
            when "10110111" => ctl <= "0010000000000000000000";
            when "10111000" => ctl <= "0010000000000000000000";
            when "10111001" => ctl <= "0010000000000000000000";
            when "10111010" => ctl <= "0010000000000000000000";
            when "10111011" => ctl <= "0010000000000000000000";
            when "10111100" => ctl <= "0010000000000000000000";
            when "10111101" => ctl <= "0010000000000000000000";
            when "10111110" => ctl <= "0010000000000000000000";
            when "10111111" => ctl <= "0010000000000000000000";

            when "11000000" => ctl <= "0010000000000000000000";
            when "11000001" => ctl <= "0010000000000000000000";
            when "11000010" => ctl <= "0010000000000000000000";
            when "11000011" => ctl <= "0010000000000000000000";
            when "11000100" => ctl <= "0010000000000000000000";
            when "11000101" => ctl <= "0001100110110010001001";
            when "11000110" => ctl <= "0010000000000000000000";
            when "11000111" => ctl <= "0010000000000000000000";
            when "11001000" => ctl <= "0010000000000000000000";
            when "11001001" => ctl <= "0010000000000000000000";
            when "11001010" => ctl <= "0010000000000000000000";
            when "11001011" => ctl <= "0010000000000000000000";
            when "11001100" => ctl <= "0010000000000000000000";
            when "11001101" => ctl <= "0010000000000000000000";
            when "11001110" => ctl <= "0010000000000000000000";
            when "11001111" => ctl <= "0010000000000000000000";

            when "11010000" => ctl <= "0010000000000000000000";
            when "11010001" => ctl <= "0010000000000000000000";
            when "11010010" => ctl <= "0010000000000000000000";
            when "11010011" => ctl <= "0010000000000000000000";
            when "11010100" => ctl <= "0010000000000000000000";
            when "11010101" => ctl <= "0010000000000000000000";
            when "11010110" => ctl <= "0010000000000000000000";
            when "11010111" => ctl <= "0010000000000000000000";
            when "11011000" => ctl <= "0010000000000000000000";
            when "11011001" => ctl <= "0010000000000000000000";
            when "11011010" => ctl <= "0010000000000000000000";
            when "11011011" => ctl <= "0010000000000000000000";
            when "11011100" => ctl <= "0010000000000000000000";
            when "11011101" => ctl <= "0010000000000000000000";
            when "11011110" => ctl <= "0010000000000000000000";
            when "11011111" => ctl <= "0010000000000000000000";

            when "11100000" => ctl <= "0010000000000000000000";
            when "11100001" => ctl <= "0010000000000000000000";
            when "11100010" => ctl <= "0010000000000000000000";
            when "11100011" => ctl <= "0010000000000000000000";
            when "11100100" => ctl <= "0010000000000000000000";
            when "11100101" => ctl <= "0001100111110010001001";
            when "11100110" => ctl <= "0010000000000000000000";
            when "11100111" => ctl <= "0010000000000000000000";
            when "11101000" => ctl <= "0010000000000000000000";
            when "11101001" => ctl <= "0010000000000000000000";
            when "11101010" => ctl <= "0010000000000000000000";
            when "11101011" => ctl <= "0010000000000000000000";
            when "11101100" => ctl <= "0010000000000000000000";
            when "11101101" => ctl <= "0010000000000000000000";
            when "11101110" => ctl <= "0010000000000000000000";
            when "11101111" => ctl <= "0010000000000000000000";

            when "11110000" => ctl <= "0010000000000000000000";
            when "11110001" => ctl <= "0010000000000000000000";
            when "11110010" => ctl <= "0010000000000000000000";
            when "11110011" => ctl <= "0010000000000000000000";
            when "11110100" => ctl <= "0010000000000000000000";
            when "11110101" => ctl <= "0010000000000000000000";
            when "11110110" => ctl <= "0010000000000000000000";
            when "11110111" => ctl <= "0010000000000000000000";
            when "11111000" => ctl <= "0010000000000000000000";
            when "11111001" => ctl <= "0010000000000000000000";
            when "11111010" => ctl <= "0010000000000000000000";
            when "11111011" => ctl <= "0010000000000000000000";
            when "11111100" => ctl <= "0010000000000000000000";
            when "11111101" => ctl <= "0010000000000000000000";
            when "11111110" => ctl <= "0010000000000000000000";
            when "11111111" => ctl <= "0010000000000000000000";

            -- Default to avoid latch
            when others => ctl <= "0010000000000000000000";
         end case;
      end if;

      if cnt_r = 3 then
         case inst_r is
            when "00000000" => ctl <= "0010000000000000000000";
            when "00000001" => ctl <= "0010000000000000000000";
            when "00000010" => ctl <= "0010000000000000000000";
            when "00000011" => ctl <= "0010000000000000000000";
            when "00000100" => ctl <= "0010000000000000000000";
            when "00000101" => ctl <= "0000000000000000000101";
            when "00000110" => ctl <= "0010000000000000000000";
            when "00000111" => ctl <= "0010000000000000000000";
            when "00001000" => ctl <= "0010000000000000000000";
            when "00001001" => ctl <= "0010000000000000000000";
            when "00001010" => ctl <= "0010000000000000000000";
            when "00001011" => ctl <= "0010000000000000000000";
            when "00001100" => ctl <= "0010000000000000000000";
            when "00001101" => ctl <= "0010000000000000000000";
            when "00001110" => ctl <= "0010000000000000000000";
            when "00001111" => ctl <= "0010000000000000000000";

            when "00010000" => ctl <= "0010000000000000000000";
            when "00010001" => ctl <= "0010000000000000000000";
            when "00010010" => ctl <= "0010000000000000000000";
            when "00010011" => ctl <= "0010000000000000000000";
            when "00010100" => ctl <= "0010000000000000000000";
            when "00010101" => ctl <= "0010000000000000000000";
            when "00010110" => ctl <= "0010000000000000000000";
            when "00010111" => ctl <= "0010000000000000000000";
            when "00011000" => ctl <= "0010000000000000000000";
            when "00011001" => ctl <= "0010000000000000000000";
            when "00011010" => ctl <= "0010000000000000000000";
            when "00011011" => ctl <= "0010000000000000000000";
            when "00011100" => ctl <= "0010000000000000000000";
            when "00011101" => ctl <= "0010000000000000000000";
            when "00011110" => ctl <= "0010000000000000000000";
            when "00011111" => ctl <= "0010000000000000000000";

            when "00100000" => ctl <= "0010000000000000000000";
            when "00100001" => ctl <= "0010000000000000000000";
            when "00100010" => ctl <= "0010000000000000000000";
            when "00100011" => ctl <= "0010000000000000000000";
            when "00100100" => ctl <= "0010000000000000000000";
            when "00100101" => ctl <= "0000000000000000000101";
            when "00100110" => ctl <= "0010000000000000000000";
            when "00100111" => ctl <= "0010000000000000000000";
            when "00101000" => ctl <= "0010000000000000000000";
            when "00101001" => ctl <= "0010000000000000000000";
            when "00101010" => ctl <= "0010000000000000000000";
            when "00101011" => ctl <= "0010000000000000000000";
            when "00101100" => ctl <= "0010000000000000000000";
            when "00101101" => ctl <= "0010000000000000000000";
            when "00101110" => ctl <= "0010000000000000000000";
            when "00101111" => ctl <= "0010000000000000000000";

            when "00110000" => ctl <= "0010000000000000000000";
            when "00110001" => ctl <= "0010000000000000000000";
            when "00110010" => ctl <= "0010000000000000000000";
            when "00110011" => ctl <= "0010000000000000000000";
            when "00110100" => ctl <= "0010000000000000000000";
            when "00110101" => ctl <= "0010000000000000000000";
            when "00110110" => ctl <= "0010000000000000000000";
            when "00110111" => ctl <= "0010000000000000000000";
            when "00111000" => ctl <= "0010000000000000000000";
            when "00111001" => ctl <= "0010000000000000000000";
            when "00111010" => ctl <= "0010000000000000000000";
            when "00111011" => ctl <= "0010000000000000000000";
            when "00111100" => ctl <= "0010000000000000000000";
            when "00111101" => ctl <= "0010000000000000000000";
            when "00111110" => ctl <= "0010000000000000000000";
            when "00111111" => ctl <= "0010000000000000000000";

            when "01000000" => ctl <= "0010000000000000000000";
            when "01000001" => ctl <= "0010000000000000000000";
            when "01000010" => ctl <= "0010000000000000000000";
            when "01000011" => ctl <= "0010000000000000000000";
            when "01000100" => ctl <= "0010000000000000000000";
            when "01000101" => ctl <= "0000000000000000000101";
            when "01000110" => ctl <= "0010000000000000000000";
            when "01000111" => ctl <= "0010000000000000000000";
            when "01001000" => ctl <= "0010000000000000000000";
            when "01001001" => ctl <= "0010000000000000000000";
            when "01001010" => ctl <= "0010000000000000000000";
            when "01001011" => ctl <= "0010000000000000000000";
            when "01001100" => ctl <= "0010000000000000000000";
            when "01001101" => ctl <= "0010000000000000000000";
            when "01001110" => ctl <= "0010000000000000000000";
            when "01001111" => ctl <= "0010000000000000000000";

            when "01010000" => ctl <= "0010000000000000000000";
            when "01010001" => ctl <= "0010000000000000000000";
            when "01010010" => ctl <= "0010000000000000000000";
            when "01010011" => ctl <= "0010000000000000000000";
            when "01010100" => ctl <= "0010000000000000000000";
            when "01010101" => ctl <= "0010000000000000000000";
            when "01010110" => ctl <= "0010000000000000000000";
            when "01010111" => ctl <= "0010000000000000000000";
            when "01011000" => ctl <= "0010000000000000000000";
            when "01011001" => ctl <= "0010000000000000000000";
            when "01011010" => ctl <= "0010000000000000000000";
            when "01011011" => ctl <= "0010000000000000000000";
            when "01011100" => ctl <= "0010000000000000000000";
            when "01011101" => ctl <= "0010000000000000000000";
            when "01011110" => ctl <= "0010000000000000000000";
            when "01011111" => ctl <= "0010000000000000000000";

            when "01100000" => ctl <= "0010000000000000000000";
            when "01100001" => ctl <= "0010000000000000000000";
            when "01100010" => ctl <= "0010000000000000000000";
            when "01100011" => ctl <= "0010000000000000000000";
            when "01100100" => ctl <= "0010000000000000000000";
            when "01100101" => ctl <= "0000000000000000000101";
            when "01100110" => ctl <= "0010000000000000000000";
            when "01100111" => ctl <= "0010000000000000000000";
            when "01101000" => ctl <= "0010000000000000000000";
            when "01101001" => ctl <= "0010000000000000000000";
            when "01101010" => ctl <= "0010000000000000000000";
            when "01101011" => ctl <= "0010000000000000000000";
            when "01101100" => ctl <= "0010000000000000000000";
            when "01101101" => ctl <= "0010000000000000000000";
            when "01101110" => ctl <= "0010000000000000000000";
            when "01101111" => ctl <= "0010000000000000000000";

            when "01110000" => ctl <= "0010000000000000000000";
            when "01110001" => ctl <= "0010000000000000000000";
            when "01110010" => ctl <= "0010000000000000000000";
            when "01110011" => ctl <= "0010000000000000000000";
            when "01110100" => ctl <= "0010000000000000000000";
            when "01110101" => ctl <= "0010000000000000000000";
            when "01110110" => ctl <= "0010000000000000000000";
            when "01110111" => ctl <= "0010000000000000000000";
            when "01111000" => ctl <= "0010000000000000000000";
            when "01111001" => ctl <= "0010000000000000000000";
            when "01111010" => ctl <= "0010000000000000000000";
            when "01111011" => ctl <= "0010000000000000000000";
            when "01111100" => ctl <= "0010000000000000000000";
            when "01111101" => ctl <= "0010000000000000000000";
            when "01111110" => ctl <= "0010000000000000000000";
            when "01111111" => ctl <= "0010000000000000000000";

            when "10000000" => ctl <= "0010000000000000000000";
            when "10000001" => ctl <= "0010000000000000000000";
            when "10000010" => ctl <= "0010000000000000000000";
            when "10000011" => ctl <= "0010000000000000000000";
            when "10000100" => ctl <= "0010000000000000000000";
            when "10000101" => ctl <= "0000000000000000000110";
            when "10000110" => ctl <= "0010000000000000000000";
            when "10000111" => ctl <= "0010000000000000000000";
            when "10001000" => ctl <= "0010000000000000000000";
            when "10001001" => ctl <= "0010000000000000000000";
            when "10001010" => ctl <= "0010000000000000000000";
            when "10001011" => ctl <= "0010000000000000000000";
            when "10001100" => ctl <= "0010000000000000000000";
            when "10001101" => ctl <= "0010000000000000000000";
            when "10001110" => ctl <= "0010000000000000000000";
            when "10001111" => ctl <= "0010000000000000000000";

            when "10010000" => ctl <= "0010000000000000000000";
            when "10010001" => ctl <= "0010000000000000000000";
            when "10010010" => ctl <= "0010000000000000000000";
            when "10010011" => ctl <= "0010000000000000000000";
            when "10010100" => ctl <= "0010000000000000000000";
            when "10010101" => ctl <= "0010000000000000000000";
            when "10010110" => ctl <= "0010000000000000000000";
            when "10010111" => ctl <= "0010000000000000000000";
            when "10011000" => ctl <= "0010000000000000000000";
            when "10011001" => ctl <= "0010000000000000000000";
            when "10011010" => ctl <= "0010000000000000000000";
            when "10011011" => ctl <= "0010000000000000000000";
            when "10011100" => ctl <= "0010000000000000000000";
            when "10011101" => ctl <= "0010000000000000000000";
            when "10011110" => ctl <= "0010000000000000000000";
            when "10011111" => ctl <= "0010000000000000000000";

            when "10100000" => ctl <= "0010000000000000000000";
            when "10100001" => ctl <= "0010000000000000000000";
            when "10100010" => ctl <= "0010000000000000000000";
            when "10100011" => ctl <= "0010000000000000000000";
            when "10100100" => ctl <= "0010000000000000000000";
            when "10100101" => ctl <= "0000000000000000000101";
            when "10100110" => ctl <= "0010000000000000000000";
            when "10100111" => ctl <= "0010000000000000000000";
            when "10101000" => ctl <= "0010000000000000000000";
            when "10101001" => ctl <= "0010000000000000000000";
            when "10101010" => ctl <= "0010000000000000000000";
            when "10101011" => ctl <= "0010000000000000000000";
            when "10101100" => ctl <= "0010000000000000000000";
            when "10101101" => ctl <= "0010000000000000000000";
            when "10101110" => ctl <= "0010000000000000000000";
            when "10101111" => ctl <= "0010000000000000000000";

            when "10110000" => ctl <= "0010000000000000000000";
            when "10110001" => ctl <= "0010000000000000000000";
            when "10110010" => ctl <= "0010000000000000000000";
            when "10110011" => ctl <= "0010000000000000000000";
            when "10110100" => ctl <= "0010000000000000000000";
            when "10110101" => ctl <= "0010000000000000000000";
            when "10110110" => ctl <= "0010000000000000000000";
            when "10110111" => ctl <= "0010000000000000000000";
            when "10111000" => ctl <= "0010000000000000000000";
            when "10111001" => ctl <= "0010000000000000000000";
            when "10111010" => ctl <= "0010000000000000000000";
            when "10111011" => ctl <= "0010000000000000000000";
            when "10111100" => ctl <= "0010000000000000000000";
            when "10111101" => ctl <= "0010000000000000000000";
            when "10111110" => ctl <= "0010000000000000000000";
            when "10111111" => ctl <= "0010000000000000000000";

            when "11000000" => ctl <= "0010000000000000000000";
            when "11000001" => ctl <= "0010000000000000000000";
            when "11000010" => ctl <= "0010000000000000000000";
            when "11000011" => ctl <= "0010000000000000000000";
            when "11000100" => ctl <= "0010000000000000000000";
            when "11000101" => ctl <= "0000000000000000000101";
            when "11000110" => ctl <= "0010000000000000000000";
            when "11000111" => ctl <= "0010000000000000000000";
            when "11001000" => ctl <= "0010000000000000000000";
            when "11001001" => ctl <= "0010000000000000000000";
            when "11001010" => ctl <= "0010000000000000000000";
            when "11001011" => ctl <= "0010000000000000000000";
            when "11001100" => ctl <= "0010000000000000000000";
            when "11001101" => ctl <= "0010000000000000000000";
            when "11001110" => ctl <= "0010000000000000000000";
            when "11001111" => ctl <= "0010000000000000000000";

            when "11010000" => ctl <= "0010000000000000000000";
            when "11010001" => ctl <= "0010000000000000000000";
            when "11010010" => ctl <= "0010000000000000000000";
            when "11010011" => ctl <= "0010000000000000000000";
            when "11010100" => ctl <= "0010000000000000000000";
            when "11010101" => ctl <= "0010000000000000000000";
            when "11010110" => ctl <= "0010000000000000000000";
            when "11010111" => ctl <= "0010000000000000000000";
            when "11011000" => ctl <= "0010000000000000000000";
            when "11011001" => ctl <= "0010000000000000000000";
            when "11011010" => ctl <= "0010000000000000000000";
            when "11011011" => ctl <= "0010000000000000000000";
            when "11011100" => ctl <= "0010000000000000000000";
            when "11011101" => ctl <= "0010000000000000000000";
            when "11011110" => ctl <= "0010000000000000000000";
            when "11011111" => ctl <= "0010000000000000000000";

            when "11100000" => ctl <= "0010000000000000000000";
            when "11100001" => ctl <= "0010000000000000000000";
            when "11100010" => ctl <= "0010000000000000000000";
            when "11100011" => ctl <= "0010000000000000000000";
            when "11100100" => ctl <= "0010000000000000000000";
            when "11100101" => ctl <= "0000000000000000000101";
            when "11100110" => ctl <= "0010000000000000000000";
            when "11100111" => ctl <= "0010000000000000000000";
            when "11101000" => ctl <= "0010000000000000000000";
            when "11101001" => ctl <= "0010000000000000000000";
            when "11101010" => ctl <= "0010000000000000000000";
            when "11101011" => ctl <= "0010000000000000000000";
            when "11101100" => ctl <= "0010000000000000000000";
            when "11101101" => ctl <= "0010000000000000000000";
            when "11101110" => ctl <= "0010000000000000000000";
            when "11101111" => ctl <= "0010000000000000000000";

            when "11110000" => ctl <= "0010000000000000000000";
            when "11110001" => ctl <= "0010000000000000000000";
            when "11110010" => ctl <= "0010000000000000000000";
            when "11110011" => ctl <= "0010000000000000000000";
            when "11110100" => ctl <= "0010000000000000000000";
            when "11110101" => ctl <= "0010000000000000000000";
            when "11110110" => ctl <= "0010000000000000000000";
            when "11110111" => ctl <= "0010000000000000000000";
            when "11111000" => ctl <= "0010000000000000000000";
            when "11111001" => ctl <= "0010000000000000000000";
            when "11111010" => ctl <= "0010000000000000000000";
            when "11111011" => ctl <= "0010000000000000000000";
            when "11111100" => ctl <= "0010000000000000000000";
            when "11111101" => ctl <= "0010000000000000000000";
            when "11111110" => ctl <= "0010000000000000000000";
            when "11111111" => ctl <= "0010000000000000000000";

            -- Default to avoid latch
            when others     => ctl <= "0010000000000000000000";
         end case;
      end if;

      if cnt_r = 4 then
         case inst_r is
            when "00000000" => ctl <= "0010000000000000000000";
            when "00000001" => ctl <= "0010000000000000000000";
            when "00000010" => ctl <= "0010000000000000000000";
            when "00000011" => ctl <= "0010000000000000000000";
            when "00000100" => ctl <= "0010000000000000000000";
            when "00000101" => ctl <= "0000000000000000000101";
            when "00000110" => ctl <= "0010000000000000000000";
            when "00000111" => ctl <= "0010000000000000000000";
            when "00001000" => ctl <= "0010000000000000000000";
            when "00001001" => ctl <= "0010000000000000000000";
            when "00001010" => ctl <= "0010000000000000000000";
            when "00001011" => ctl <= "0010000000000000000000";
            when "00001100" => ctl <= "0010000000000000000000";
            when "00001101" => ctl <= "0010000000000000000000";
            when "00001110" => ctl <= "0010000000000000000000";
            when "00001111" => ctl <= "0010000000000000000000";

            when "00010000" => ctl <= "0010000000000000000000";
            when "00010001" => ctl <= "0010000000000000000000";
            when "00010010" => ctl <= "0010000000000000000000";
            when "00010011" => ctl <= "0010000000000000000000";
            when "00010100" => ctl <= "0010000000000000000000";
            when "00010101" => ctl <= "0010000000000000000000";
            when "00010110" => ctl <= "0010000000000000000000";
            when "00010111" => ctl <= "0010000000000000000000";
            when "00011000" => ctl <= "0010000000000000000000";
            when "00011001" => ctl <= "0010000000000000000000";
            when "00011010" => ctl <= "0010000000000000000000";
            when "00011011" => ctl <= "0010000000000000000000";
            when "00011100" => ctl <= "0010000000000000000000";
            when "00011101" => ctl <= "0010000000000000000000";
            when "00011110" => ctl <= "0010000000000000000000";
            when "00011111" => ctl <= "0010000000000000000000";

            when "00100000" => ctl <= "0010000000000000000000";
            when "00100001" => ctl <= "0010000000000000000000";
            when "00100010" => ctl <= "0010000000000000000000";
            when "00100011" => ctl <= "0010000000000000000000";
            when "00100100" => ctl <= "0010000000000000000000";
            when "00100101" => ctl <= "0000000000000000000101";
            when "00100110" => ctl <= "0010000000000000000000";
            when "00100111" => ctl <= "0010000000000000000000";
            when "00101000" => ctl <= "0010000000000000000000";
            when "00101001" => ctl <= "0010000000000000000000";
            when "00101010" => ctl <= "0010000000000000000000";
            when "00101011" => ctl <= "0010000000000000000000";
            when "00101100" => ctl <= "0010000000000000000000";
            when "00101101" => ctl <= "0010000000000000000000";
            when "00101110" => ctl <= "0010000000000000000000";
            when "00101111" => ctl <= "0010000000000000000000";

            when "00110000" => ctl <= "0010000000000000000000";
            when "00110001" => ctl <= "0010000000000000000000";
            when "00110010" => ctl <= "0010000000000000000000";
            when "00110011" => ctl <= "0010000000000000000000";
            when "00110100" => ctl <= "0010000000000000000000";
            when "00110101" => ctl <= "0010000000000000000000";
            when "00110110" => ctl <= "0010000000000000000000";
            when "00110111" => ctl <= "0010000000000000000000";
            when "00111000" => ctl <= "0010000000000000000000";
            when "00111001" => ctl <= "0010000000000000000000";
            when "00111010" => ctl <= "0010000000000000000000";
            when "00111011" => ctl <= "0010000000000000000000";
            when "00111100" => ctl <= "0010000000000000000000";
            when "00111101" => ctl <= "0010000000000000000000";
            when "00111110" => ctl <= "0010000000000000000000";
            when "00111111" => ctl <= "0010000000000000000000";

            when "01000000" => ctl <= "0010000000000000000000";
            when "01000001" => ctl <= "0010000000000000000000";
            when "01000010" => ctl <= "0010000000000000000000";
            when "01000011" => ctl <= "0010000000000000000000";
            when "01000100" => ctl <= "0010000000000000000000";
            when "01000101" => ctl <= "0000000000000000000101";
            when "01000110" => ctl <= "0010000000000000000000";
            when "01000111" => ctl <= "0010000000000000000000";
            when "01001000" => ctl <= "0010000000000000000000";
            when "01001001" => ctl <= "0010000000000000000000";
            when "01001010" => ctl <= "0010000000000000000000";
            when "01001011" => ctl <= "0010000000000000000000";
            when "01001100" => ctl <= "0010000000000000000000";
            when "01001101" => ctl <= "0010000000000000000000";
            when "01001110" => ctl <= "0010000000000000000000";
            when "01001111" => ctl <= "0010000000000000000000";

            when "01010000" => ctl <= "0010000000000000000000";
            when "01010001" => ctl <= "0010000000000000000000";
            when "01010010" => ctl <= "0010000000000000000000";
            when "01010011" => ctl <= "0010000000000000000000";
            when "01010100" => ctl <= "0010000000000000000000";
            when "01010101" => ctl <= "0010000000000000000000";
            when "01010110" => ctl <= "0010000000000000000000";
            when "01010111" => ctl <= "0010000000000000000000";
            when "01011000" => ctl <= "0010000000000000000000";
            when "01011001" => ctl <= "0010000000000000000000";
            when "01011010" => ctl <= "0010000000000000000000";
            when "01011011" => ctl <= "0010000000000000000000";
            when "01011100" => ctl <= "0010000000000000000000";
            when "01011101" => ctl <= "0010000000000000000000";
            when "01011110" => ctl <= "0010000000000000000000";
            when "01011111" => ctl <= "0010000000000000000000";

            when "01100000" => ctl <= "0010000000000000000000";
            when "01100001" => ctl <= "0010000000000000000000";
            when "01100010" => ctl <= "0010000000000000000000";
            when "01100011" => ctl <= "0010000000000000000000";
            when "01100100" => ctl <= "0010000000000000000000";
            when "01100101" => ctl <= "0000000000000000000101";
            when "01100110" => ctl <= "0010000000000000000000";
            when "01100111" => ctl <= "0010000000000000000000";
            when "01101000" => ctl <= "0010000000000000000000";
            when "01101001" => ctl <= "0010000000000000000000";
            when "01101010" => ctl <= "0010000000000000000000";
            when "01101011" => ctl <= "0010000000000000000000";
            when "01101100" => ctl <= "0010000000000000000000";
            when "01101101" => ctl <= "0010000000000000000000";
            when "01101110" => ctl <= "0010000000000000000000";
            when "01101111" => ctl <= "0010000000000000000000";

            when "01110000" => ctl <= "0010000000000000000000";
            when "01110001" => ctl <= "0010000000000000000000";
            when "01110010" => ctl <= "0010000000000000000000";
            when "01110011" => ctl <= "0010000000000000000000";
            when "01110100" => ctl <= "0010000000000000000000";
            when "01110101" => ctl <= "0010000000000000000000";
            when "01110110" => ctl <= "0010000000000000000000";
            when "01110111" => ctl <= "0010000000000000000000";
            when "01111000" => ctl <= "0010000000000000000000";
            when "01111001" => ctl <= "0010000000000000000000";
            when "01111010" => ctl <= "0010000000000000000000";
            when "01111011" => ctl <= "0010000000000000000000";
            when "01111100" => ctl <= "0010000000000000000000";
            when "01111101" => ctl <= "0010000000000000000000";
            when "01111110" => ctl <= "0010000000000000000000";
            when "01111111" => ctl <= "0010000000000000000000";

            when "10000000" => ctl <= "0010000000000000000000";
            when "10000001" => ctl <= "0010000000000000000000";
            when "10000010" => ctl <= "0010000000000000000000";
            when "10000011" => ctl <= "0010000000000000000000";
            when "10000100" => ctl <= "0010000000000000000000";
            when "10000101" => ctl <= "0000000000000000000110";
            when "10000110" => ctl <= "0010000000000000000000";
            when "10000111" => ctl <= "0010000000000000000000";
            when "10001000" => ctl <= "0010000000000000000000";
            when "10001001" => ctl <= "0010000000000000000000";
            when "10001010" => ctl <= "0010000000000000000000";
            when "10001011" => ctl <= "0010000000000000000000";
            when "10001100" => ctl <= "0010000000000000000000";
            when "10001101" => ctl <= "0010000000000000000000";
            when "10001110" => ctl <= "0010000000000000000000";
            when "10001111" => ctl <= "0010000000000000000000";

            when "10010000" => ctl <= "0010000000000000000000";
            when "10010001" => ctl <= "0010000000000000000000";
            when "10010010" => ctl <= "0010000000000000000000";
            when "10010011" => ctl <= "0010000000000000000000";
            when "10010100" => ctl <= "0010000000000000000000";
            when "10010101" => ctl <= "0010000000000000000000";
            when "10010110" => ctl <= "0010000000000000000000";
            when "10010111" => ctl <= "0010000000000000000000";
            when "10011000" => ctl <= "0010000000000000000000";
            when "10011001" => ctl <= "0010000000000000000000";
            when "10011010" => ctl <= "0010000000000000000000";
            when "10011011" => ctl <= "0010000000000000000000";
            when "10011100" => ctl <= "0010000000000000000000";
            when "10011101" => ctl <= "0010000000000000000000";
            when "10011110" => ctl <= "0010000000000000000000";
            when "10011111" => ctl <= "0010000000000000000000";

            when "10100000" => ctl <= "0010000000000000000000";
            when "10100001" => ctl <= "0010000000000000000000";
            when "10100010" => ctl <= "0010000000000000000000";
            when "10100011" => ctl <= "0010000000000000000000";
            when "10100100" => ctl <= "0010000000000000000000";
            when "10100101" => ctl <= "0000000000000000000101";
            when "10100110" => ctl <= "0010000000000000000000";
            when "10100111" => ctl <= "0010000000000000000000";
            when "10101000" => ctl <= "0010000000000000000000";
            when "10101001" => ctl <= "0010000000000000000000";
            when "10101010" => ctl <= "0010000000000000000000";
            when "10101011" => ctl <= "0010000000000000000000";
            when "10101100" => ctl <= "0010000000000000000000";
            when "10101101" => ctl <= "0010000000000000000000";
            when "10101110" => ctl <= "0010000000000000000000";
            when "10101111" => ctl <= "0010000000000000000000";

            when "10110000" => ctl <= "0010000000000000000000";
            when "10110001" => ctl <= "0010000000000000000000";
            when "10110010" => ctl <= "0010000000000000000000";
            when "10110011" => ctl <= "0010000000000000000000";
            when "10110100" => ctl <= "0010000000000000000000";
            when "10110101" => ctl <= "0010000000000000000000";
            when "10110110" => ctl <= "0010000000000000000000";
            when "10110111" => ctl <= "0010000000000000000000";
            when "10111000" => ctl <= "0010000000000000000000";
            when "10111001" => ctl <= "0010000000000000000000";
            when "10111010" => ctl <= "0010000000000000000000";
            when "10111011" => ctl <= "0010000000000000000000";
            when "10111100" => ctl <= "0010000000000000000000";
            when "10111101" => ctl <= "0010000000000000000000";
            when "10111110" => ctl <= "0010000000000000000000";
            when "10111111" => ctl <= "0010000000000000000000";

            when "11000000" => ctl <= "0010000000000000000000";
            when "11000001" => ctl <= "0010000000000000000000";
            when "11000010" => ctl <= "0010000000000000000000";
            when "11000011" => ctl <= "0010000000000000000000";
            when "11000100" => ctl <= "0010000000000000000000";
            when "11000101" => ctl <= "0000000000000000000101";
            when "11000110" => ctl <= "0010000000000000000000";
            when "11000111" => ctl <= "0010000000000000000000";
            when "11001000" => ctl <= "0010000000000000000000";
            when "11001001" => ctl <= "0010000000000000000000";
            when "11001010" => ctl <= "0010000000000000000000";
            when "11001011" => ctl <= "0010000000000000000000";
            when "11001100" => ctl <= "0010000000000000000000";
            when "11001101" => ctl <= "0010000000000000000000";
            when "11001110" => ctl <= "0010000000000000000000";
            when "11001111" => ctl <= "0010000000000000000000";

            when "11010000" => ctl <= "0010000000000000000000";
            when "11010001" => ctl <= "0010000000000000000000";
            when "11010010" => ctl <= "0010000000000000000000";
            when "11010011" => ctl <= "0010000000000000000000";
            when "11010100" => ctl <= "0010000000000000000000";
            when "11010101" => ctl <= "0010000000000000000000";
            when "11010110" => ctl <= "0010000000000000000000";
            when "11010111" => ctl <= "0010000000000000000000";
            when "11011000" => ctl <= "0010000000000000000000";
            when "11011001" => ctl <= "0010000000000000000000";
            when "11011010" => ctl <= "0010000000000000000000";
            when "11011011" => ctl <= "0010000000000000000000";
            when "11011100" => ctl <= "0010000000000000000000";
            when "11011101" => ctl <= "0010000000000000000000";
            when "11011110" => ctl <= "0010000000000000000000";
            when "11011111" => ctl <= "0010000000000000000000";

            when "11100000" => ctl <= "0010000000000000000000";
            when "11100001" => ctl <= "0010000000000000000000";
            when "11100010" => ctl <= "0010000000000000000000";
            when "11100011" => ctl <= "0010000000000000000000";
            when "11100100" => ctl <= "0010000000000000000000";
            when "11100101" => ctl <= "0000000000000000000101";
            when "11100110" => ctl <= "0010000000000000000000";
            when "11100111" => ctl <= "0010000000000000000000";
            when "11101000" => ctl <= "0010000000000000000000";
            when "11101001" => ctl <= "0010000000000000000000";
            when "11101010" => ctl <= "0010000000000000000000";
            when "11101011" => ctl <= "0010000000000000000000";
            when "11101100" => ctl <= "0010000000000000000000";
            when "11101101" => ctl <= "0010000000000000000000";
            when "11101110" => ctl <= "0010000000000000000000";
            when "11101111" => ctl <= "0010000000000000000000";

            when "11110000" => ctl <= "0010000000000000000000";
            when "11110001" => ctl <= "0010000000000000000000";
            when "11110010" => ctl <= "0010000000000000000000";
            when "11110011" => ctl <= "0010000000000000000000";
            when "11110100" => ctl <= "0010000000000000000000";
            when "11110101" => ctl <= "0010000000000000000000";
            when "11110110" => ctl <= "0010000000000000000000";
            when "11110111" => ctl <= "0010000000000000000000";
            when "11111000" => ctl <= "0010000000000000000000";
            when "11111001" => ctl <= "0010000000000000000000";
            when "11111010" => ctl <= "0010000000000000000000";
            when "11111011" => ctl <= "0010000000000000000000";
            when "11111100" => ctl <= "0010000000000000000000";
            when "11111101" => ctl <= "0010000000000000000000";
            when "11111110" => ctl <= "0010000000000000000000";
            when "11111111" => ctl <= "0010000000000000000000";

            -- Default to avoid latch
            when others     => ctl <= "0010000000000000000000";
         end case;
      end if;

      if cnt_r = 5 then
         case inst_r is
            when "00000000" => ctl <= "0010000000000000000000";
            when "00000001" => ctl <= "0010000000000000000000";
            when "00000010" => ctl <= "0010000000000000000000";
            when "00000011" => ctl <= "0010000000000000000000";
            when "00000100" => ctl <= "0010000000000000000000";
            when "00000101" => ctl <= "0000000000000000000101";
            when "00000110" => ctl <= "0010000000000000000000";
            when "00000111" => ctl <= "0010000000000000000000";
            when "00001000" => ctl <= "0010000000000000000000";
            when "00001001" => ctl <= "0010000000000000000000";
            when "00001010" => ctl <= "0010000000000000000000";
            when "00001011" => ctl <= "0010000000000000000000";
            when "00001100" => ctl <= "0010000000000000000000";
            when "00001101" => ctl <= "0010000000000000000000";
            when "00001110" => ctl <= "0010000000000000000000";
            when "00001111" => ctl <= "0010000000000000000000";

            when "00010000" => ctl <= "0010000000000000000000";
            when "00010001" => ctl <= "0010000000000000000000";
            when "00010010" => ctl <= "0010000000000000000000";
            when "00010011" => ctl <= "0010000000000000000000";
            when "00010100" => ctl <= "0010000000000000000000";
            when "00010101" => ctl <= "0010000000000000000000";
            when "00010110" => ctl <= "0010000000000000000000";
            when "00010111" => ctl <= "0010000000000000000000";
            when "00011000" => ctl <= "0010000000000000000000";
            when "00011001" => ctl <= "0010000000000000000000";
            when "00011010" => ctl <= "0010000000000000000000";
            when "00011011" => ctl <= "0010000000000000000000";
            when "00011100" => ctl <= "0010000000000000000000";
            when "00011101" => ctl <= "0010000000000000000000";
            when "00011110" => ctl <= "0010000000000000000000";
            when "00011111" => ctl <= "0010000000000000000000";

            when "00100000" => ctl <= "0010000000000000000000";
            when "00100001" => ctl <= "0010000000000000000000";
            when "00100010" => ctl <= "0010000000000000000000";
            when "00100011" => ctl <= "0010000000000000000000";
            when "00100100" => ctl <= "0010000000000000000000";
            when "00100101" => ctl <= "0000000000000000000101";
            when "00100110" => ctl <= "0010000000000000000000";
            when "00100111" => ctl <= "0010000000000000000000";
            when "00101000" => ctl <= "0010000000000000000000";
            when "00101001" => ctl <= "0010000000000000000000";
            when "00101010" => ctl <= "0010000000000000000000";
            when "00101011" => ctl <= "0010000000000000000000";
            when "00101100" => ctl <= "0010000000000000000000";
            when "00101101" => ctl <= "0010000000000000000000";
            when "00101110" => ctl <= "0010000000000000000000";
            when "00101111" => ctl <= "0010000000000000000000";

            when "00110000" => ctl <= "0010000000000000000000";
            when "00110001" => ctl <= "0010000000000000000000";
            when "00110010" => ctl <= "0010000000000000000000";
            when "00110011" => ctl <= "0010000000000000000000";
            when "00110100" => ctl <= "0010000000000000000000";
            when "00110101" => ctl <= "0010000000000000000000";
            when "00110110" => ctl <= "0010000000000000000000";
            when "00110111" => ctl <= "0010000000000000000000";
            when "00111000" => ctl <= "0010000000000000000000";
            when "00111001" => ctl <= "0010000000000000000000";
            when "00111010" => ctl <= "0010000000000000000000";
            when "00111011" => ctl <= "0010000000000000000000";
            when "00111100" => ctl <= "0010000000000000000000";
            when "00111101" => ctl <= "0010000000000000000000";
            when "00111110" => ctl <= "0010000000000000000000";
            when "00111111" => ctl <= "0010000000000000000000";

            when "01000000" => ctl <= "0010000000000000000000";
            when "01000001" => ctl <= "0010000000000000000000";
            when "01000010" => ctl <= "0010000000000000000000";
            when "01000011" => ctl <= "0010000000000000000000";
            when "01000100" => ctl <= "0010000000000000000000";
            when "01000101" => ctl <= "0000000000000000000101";
            when "01000110" => ctl <= "0010000000000000000000";
            when "01000111" => ctl <= "0010000000000000000000";
            when "01001000" => ctl <= "0010000000000000000000";
            when "01001001" => ctl <= "0010000000000000000000";
            when "01001010" => ctl <= "0010000000000000000000";
            when "01001011" => ctl <= "0010000000000000000000";
            when "01001100" => ctl <= "0010000000000000000000";
            when "01001101" => ctl <= "0010000000000000000000";
            when "01001110" => ctl <= "0010000000000000000000";
            when "01001111" => ctl <= "0010000000000000000000";

            when "01010000" => ctl <= "0010000000000000000000";
            when "01010001" => ctl <= "0010000000000000000000";
            when "01010010" => ctl <= "0010000000000000000000";
            when "01010011" => ctl <= "0010000000000000000000";
            when "01010100" => ctl <= "0010000000000000000000";
            when "01010101" => ctl <= "0010000000000000000000";
            when "01010110" => ctl <= "0010000000000000000000";
            when "01010111" => ctl <= "0010000000000000000000";
            when "01011000" => ctl <= "0010000000000000000000";
            when "01011001" => ctl <= "0010000000000000000000";
            when "01011010" => ctl <= "0010000000000000000000";
            when "01011011" => ctl <= "0010000000000000000000";
            when "01011100" => ctl <= "0010000000000000000000";
            when "01011101" => ctl <= "0010000000000000000000";
            when "01011110" => ctl <= "0010000000000000000000";
            when "01011111" => ctl <= "0010000000000000000000";

            when "01100000" => ctl <= "0010000000000000000000";
            when "01100001" => ctl <= "0010000000000000000000";
            when "01100010" => ctl <= "0010000000000000000000";
            when "01100011" => ctl <= "0010000000000000000000";
            when "01100100" => ctl <= "0010000000000000000000";
            when "01100101" => ctl <= "0000000000000000000101";
            when "01100110" => ctl <= "0010000000000000000000";
            when "01100111" => ctl <= "0010000000000000000000";
            when "01101000" => ctl <= "0010000000000000000000";
            when "01101001" => ctl <= "0010000000000000000000";
            when "01101010" => ctl <= "0010000000000000000000";
            when "01101011" => ctl <= "0010000000000000000000";
            when "01101100" => ctl <= "0010000000000000000000";
            when "01101101" => ctl <= "0010000000000000000000";
            when "01101110" => ctl <= "0010000000000000000000";
            when "01101111" => ctl <= "0010000000000000000000";

            when "01110000" => ctl <= "0010000000000000000000";
            when "01110001" => ctl <= "0010000000000000000000";
            when "01110010" => ctl <= "0010000000000000000000";
            when "01110011" => ctl <= "0010000000000000000000";
            when "01110100" => ctl <= "0010000000000000000000";
            when "01110101" => ctl <= "0010000000000000000000";
            when "01110110" => ctl <= "0010000000000000000000";
            when "01110111" => ctl <= "0010000000000000000000";
            when "01111000" => ctl <= "0010000000000000000000";
            when "01111001" => ctl <= "0010000000000000000000";
            when "01111010" => ctl <= "0010000000000000000000";
            when "01111011" => ctl <= "0010000000000000000000";
            when "01111100" => ctl <= "0010000000000000000000";
            when "01111101" => ctl <= "0010000000000000000000";
            when "01111110" => ctl <= "0010000000000000000000";
            when "01111111" => ctl <= "0010000000000000000000";

            when "10000000" => ctl <= "0010000000000000000000";
            when "10000001" => ctl <= "0010000000000000000000";
            when "10000010" => ctl <= "0010000000000000000000";
            when "10000011" => ctl <= "0010000000000000000000";
            when "10000100" => ctl <= "0010000000000000000000";
            when "10000101" => ctl <= "0000000000000000000110";
            when "10000110" => ctl <= "0010000000000000000000";
            when "10000111" => ctl <= "0010000000000000000000";
            when "10001000" => ctl <= "0010000000000000000000";
            when "10001001" => ctl <= "0010000000000000000000";
            when "10001010" => ctl <= "0010000000000000000000";
            when "10001011" => ctl <= "0010000000000000000000";
            when "10001100" => ctl <= "0010000000000000000000";
            when "10001101" => ctl <= "0010000000000000000000";
            when "10001110" => ctl <= "0010000000000000000000";
            when "10001111" => ctl <= "0010000000000000000000";

            when "10010000" => ctl <= "0010000000000000000000";
            when "10010001" => ctl <= "0010000000000000000000";
            when "10010010" => ctl <= "0010000000000000000000";
            when "10010011" => ctl <= "0010000000000000000000";
            when "10010100" => ctl <= "0010000000000000000000";
            when "10010101" => ctl <= "0010000000000000000000";
            when "10010110" => ctl <= "0010000000000000000000";
            when "10010111" => ctl <= "0010000000000000000000";
            when "10011000" => ctl <= "0010000000000000000000";
            when "10011001" => ctl <= "0010000000000000000000";
            when "10011010" => ctl <= "0010000000000000000000";
            when "10011011" => ctl <= "0010000000000000000000";
            when "10011100" => ctl <= "0010000000000000000000";
            when "10011101" => ctl <= "0010000000000000000000";
            when "10011110" => ctl <= "0010000000000000000000";
            when "10011111" => ctl <= "0010000000000000000000";

            when "10100000" => ctl <= "0010000000000000000000";
            when "10100001" => ctl <= "0010000000000000000000";
            when "10100010" => ctl <= "0010000000000000000000";
            when "10100011" => ctl <= "0010000000000000000000";
            when "10100100" => ctl <= "0010000000000000000000";
            when "10100101" => ctl <= "0000000000000000000101";
            when "10100110" => ctl <= "0010000000000000000000";
            when "10100111" => ctl <= "0010000000000000000000";
            when "10101000" => ctl <= "0010000000000000000000";
            when "10101001" => ctl <= "0010000000000000000000";
            when "10101010" => ctl <= "0010000000000000000000";
            when "10101011" => ctl <= "0010000000000000000000";
            when "10101100" => ctl <= "0010000000000000000000";
            when "10101101" => ctl <= "0010000000000000000000";
            when "10101110" => ctl <= "0010000000000000000000";
            when "10101111" => ctl <= "0010000000000000000000";

            when "10110000" => ctl <= "0010000000000000000000";
            when "10110001" => ctl <= "0010000000000000000000";
            when "10110010" => ctl <= "0010000000000000000000";
            when "10110011" => ctl <= "0010000000000000000000";
            when "10110100" => ctl <= "0010000000000000000000";
            when "10110101" => ctl <= "0010000000000000000000";
            when "10110110" => ctl <= "0010000000000000000000";
            when "10110111" => ctl <= "0010000000000000000000";
            when "10111000" => ctl <= "0010000000000000000000";
            when "10111001" => ctl <= "0010000000000000000000";
            when "10111010" => ctl <= "0010000000000000000000";
            when "10111011" => ctl <= "0010000000000000000000";
            when "10111100" => ctl <= "0010000000000000000000";
            when "10111101" => ctl <= "0010000000000000000000";
            when "10111110" => ctl <= "0010000000000000000000";
            when "10111111" => ctl <= "0010000000000000000000";

            when "11000000" => ctl <= "0010000000000000000000";
            when "11000001" => ctl <= "0010000000000000000000";
            when "11000010" => ctl <= "0010000000000000000000";
            when "11000011" => ctl <= "0010000000000000000000";
            when "11000100" => ctl <= "0010000000000000000000";
            when "11000101" => ctl <= "0000000000000000000101";
            when "11000110" => ctl <= "0010000000000000000000";
            when "11000111" => ctl <= "0010000000000000000000";
            when "11001000" => ctl <= "0010000000000000000000";
            when "11001001" => ctl <= "0010000000000000000000";
            when "11001010" => ctl <= "0010000000000000000000";
            when "11001011" => ctl <= "0010000000000000000000";
            when "11001100" => ctl <= "0010000000000000000000";
            when "11001101" => ctl <= "0010000000000000000000";
            when "11001110" => ctl <= "0010000000000000000000";
            when "11001111" => ctl <= "0010000000000000000000";

            when "11010000" => ctl <= "0010000000000000000000";
            when "11010001" => ctl <= "0010000000000000000000";
            when "11010010" => ctl <= "0010000000000000000000";
            when "11010011" => ctl <= "0010000000000000000000";
            when "11010100" => ctl <= "0010000000000000000000";
            when "11010101" => ctl <= "0010000000000000000000";
            when "11010110" => ctl <= "0010000000000000000000";
            when "11010111" => ctl <= "0010000000000000000000";
            when "11011000" => ctl <= "0010000000000000000000";
            when "11011001" => ctl <= "0010000000000000000000";
            when "11011010" => ctl <= "0010000000000000000000";
            when "11011011" => ctl <= "0010000000000000000000";
            when "11011100" => ctl <= "0010000000000000000000";
            when "11011101" => ctl <= "0010000000000000000000";
            when "11011110" => ctl <= "0010000000000000000000";
            when "11011111" => ctl <= "0010000000000000000000";

            when "11100000" => ctl <= "0010000000000000000000";
            when "11100001" => ctl <= "0010000000000000000000";
            when "11100010" => ctl <= "0010000000000000000000";
            when "11100011" => ctl <= "0010000000000000000000";
            when "11100100" => ctl <= "0010000000000000000000";
            when "11100101" => ctl <= "0000000000000000000101";
            when "11100110" => ctl <= "0010000000000000000000";
            when "11100111" => ctl <= "0010000000000000000000";
            when "11101000" => ctl <= "0010000000000000000000";
            when "11101001" => ctl <= "0010000000000000000000";
            when "11101010" => ctl <= "0010000000000000000000";
            when "11101011" => ctl <= "0010000000000000000000";
            when "11101100" => ctl <= "0010000000000000000000";
            when "11101101" => ctl <= "0010000000000000000000";
            when "11101110" => ctl <= "0010000000000000000000";
            when "11101111" => ctl <= "0010000000000000000000";

            when "11110000" => ctl <= "0010000000000000000000";
            when "11110001" => ctl <= "0010000000000000000000";
            when "11110010" => ctl <= "0010000000000000000000";
            when "11110011" => ctl <= "0010000000000000000000";
            when "11110100" => ctl <= "0010000000000000000000";
            when "11110101" => ctl <= "0010000000000000000000";
            when "11110110" => ctl <= "0010000000000000000000";
            when "11110111" => ctl <= "0010000000000000000000";
            when "11111000" => ctl <= "0010000000000000000000";
            when "11111001" => ctl <= "0010000000000000000000";
            when "11111010" => ctl <= "0010000000000000000000";
            when "11111011" => ctl <= "0010000000000000000000";
            when "11111100" => ctl <= "0010000000000000000000";
            when "11111101" => ctl <= "0010000000000000000000";
            when "11111110" => ctl <= "0010000000000000000000";
            when "11111111" => ctl <= "0010000000000000000000";

            -- Default to avoid latch
            when others     => ctl <= "0010000000000000000000";
         end case;
      end if;
   end process;

end architecture Structural;


------------------------------------------------------------------------
-- vga_controller_640_60.vhd
------------------------------------------------------------------------
-- Author : Ulrich Zolt�n
--          Copyright 2006 Digilent, Inc.
------------------------------------------------------------------------
-- This file contains the logic to generate the synchronization signals,
-- horizontal and vertical pixel counter and video disable signal
-- for the 640x480@60Hz resolution.
------------------------------------------------------------------------
--  Behavioral description
------------------------------------------------------------------------
-- Please read the following article on the web regarding the
-- vga video timings:
-- http://www.epanorama.net/documents/pc/vga_timing.html

-- This module generates the video synch pulses for the monitor to
-- enter 640x480@60Hz resolution state. It also provides horizontal
-- and vertical counters for the currently displayed pixel and a blank
-- signal that is active when the pixel is not inside the visible screen
-- and the color outputs should be reset to 0.

-- timing diagram for the horizontal synch signal (HS)
-- 0                         648    744           800 (pixels)
-- -------------------------|______|-----------------
-- timing diagram for the vertical synch signal (VS)
-- 0                                  482    484  525 (lines)
-- -----------------------------------|______|-------

-- The blank signal is delayed one pixel clock period (40ns) from where
-- the pixel leaves the visible screen, according to the counters, to
-- account for the pixel pipeline delay. This delay happens because
-- it takes time from when the counters indicate current pixel should
-- be displayed to when the color data actually arrives at the monitor
-- pins (memory read delays, synchronization delays).
------------------------------------------------------------------------
--  Port definitions
------------------------------------------------------------------------
-- rst               - global reset signal
-- pixel_clk         - input pin, from dcm_25MHz
--                   - the clock signal generated by a DCM that has
--                   - a frequency of 25MHz.
-- HS                - output pin, to monitor
--                   - horizontal synch pulse
-- VS                - output pin, to monitor
--                   - vertical synch pulse
-- hcount            - output pin, 11 bits, to clients
--                   - horizontal count of the currently displayed
--                   - pixel (even if not in visible area)
-- vcount            - output pin, 11 bits, to clients
--                   - vertical count of the currently active video
--                   - line (even if not in visible area)
-- blank             - output pin, to clients
--                   - active when pixel is not in visible area.
------------------------------------------------------------------------
-- Revision History:
-- 09/18/2006(UlrichZ): created
------------------------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

-- the vga_ctrl entity declaration
-- read above for behavioral description and port definitions.
entity vga_ctrl is
   port(
      rst_i    : in std_logic;
      clk_i    : in std_logic;

      hs_o     : out std_logic;
      vs_o     : out std_logic;
      hcount_o : out std_logic_vector(10 downto 0);
      vcount_o : out std_logic_vector(10 downto 0);
      blank_o  : out std_logic
   );
end vga_ctrl;

architecture Behavioral of vga_ctrl is

------------------------------------------------------------------------
-- CONSTANTS
------------------------------------------------------------------------

   -- maximum value for the horizontal pixel counter
   constant HMAX  : std_logic_vector(10 downto 0) := "01100100000"; -- 800
   -- maximum value for the vertical pixel counter
   constant VMAX  : std_logic_vector(10 downto 0) := "01000001101"; -- 525
   -- total number of visible columns
   constant HLINES: std_logic_vector(10 downto 0) := "01010000000"; -- 640
   -- value for the horizontal counter where front porch ends
   constant HFP   : std_logic_vector(10 downto 0) := "01010001000"; -- 648
   -- value for the horizontal counter where the synch pulse ends
   constant HSP   : std_logic_vector(10 downto 0) := "01011101000"; -- 744
   -- total number of visible lines
   constant VLINES: std_logic_vector(10 downto 0) := "00111100000"; -- 480
   -- value for the vertical counter where the front porch ends
   constant VFP   : std_logic_vector(10 downto 0) := "00111100010"; -- 482
   -- value for the vertical counter where the synch pulse ends
   constant VSP   : std_logic_vector(10 downto 0) := "00111100100"; -- 484

   ------------------------------------------------------------------------
   -- SIGNALS
   ------------------------------------------------------------------------

   -- horizontal and vertical counters
   signal hcounter : std_logic_vector(10 downto 0) := (others => '0');
   signal vcounter : std_logic_vector(10 downto 0) := (others => '0');

   signal hs     : std_logic;
   signal vs     : std_logic;
   signal blank  : std_logic;

begin

   -- increment horizontal counter at pixel_clk rate
   -- until HMAX is reached, then reset and keep counting
   h_count: process (clk_i)
   begin
      if (rising_edge(clk_i)) then
         if (hcounter = HMAX-1) then
            hcounter <= (others => '0');
         else
            hcounter <= hcounter + 1;
         end if;

         if (rst_i = '1') then
            hcounter <= (others => '0');
         end if;
      end if;
   end process h_count;

   -- increment vertical counter when one line is finished
   -- (horizontal counter reached HMAX)
   -- until VMAX is reached, then reset and keep counting
   v_count: process(clk_i)
   begin
      if (rising_edge(clk_i)) then
         if (hcounter = HMAX-1) then
            if (vcounter = VMAX-1) then
               vcounter <= (others => '0');
            else
               vcounter <= vcounter + 1;
            end if;
         end if;

         if (rst_i = '1') then
            vcounter <= (others => '0');
         end if;
      end if;
   end process v_count;

   -- generate horizontal synch pulse
   -- when horizontal counter is between where the
   -- front porch ends and the synch pulse ends.
   -- The HS is active for a total of 96 pixels.
   hs <= '0' when (hcounter >= HFP and hcounter < HSP) 
         else '1';

   -- generate vertical synch pulse
   -- when vertical counter is between where the
   -- front porch ends and the synch pulse ends.
   -- The VS is active for a total of 2 video lines
   -- = 2*HMAX = 1600 pixels.
   vs <= '0' when (vcounter >= VFP and vcounter < VSP) 
         else '1';

   -- enable video output when pixel is in visible area
   blank <= '0' when (hcounter < HLINES and vcounter < VLINES) else '1';

   -- Register outputs
   p_output: process(clk_i)
   begin
      if(rising_edge(clk_i)) then
         hs_o     <= hs;
         vs_o     <= vs;
         hcount_o <= hcounter;
         vcount_o <= vcounter;
         blank_o  <= blank;
      end if;
   end process p_output;

end Behavioral;

library ieee;
use ieee.std_logic_1164.all;

-- This block is a dummy block that generates a number of writes from the CPU,
-- simulating the KERNAL/BASIC ROM.

entity cpu_dummy is
   port (
      clk_i     : in  std_logic;
      wr_addr_o : out std_logic_vector(2 downto 0);
      wr_en_o   : out std_logic;
      wr_data_o : out std_logic_vector(7 downto 0)
   );
end cpu_dummy;

architecture structural of cpu_dummy is

   -- This defines a type containing an array of bytes
   type wr_record is record
      addr : std_logic_vector(15 downto 0);
      data : std_logic_vector( 7 downto 0);
   end record wr_record;
   type wr_record_vector is array (natural range <>) of wr_record;

   constant wr_default : wr_record_vector := (
      -- Configure layer 1
      (X"9F25", X"00"), -- Select address port 0
      (X"9F20", X"00"),
      (X"9F21", X"30"),
      (X"9F22", X"1F"), -- Set address to 0xF3000 and increment to 1.
      (X"9F23", X"01"), -- 0xF3000
      (X"9F23", X"06"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"3E"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),

      -- Configure display composer
      (X"9F20", X"00"),
      (X"9F21", X"00"),
      (X"9F22", X"1F"), -- Set address to 0xF0000 and increment to 1.
      (X"9F23", X"01"), -- 0xF0000
      (X"9F23", X"80"),
      (X"9F23", X"80"),
      (X"9F23", X"0E"),
      (X"9F23", X"00"),
      (X"9F23", X"80"),
      (X"9F23", X"00"),
      (X"9F23", X"E0"),
      (X"9F23", X"28"),

      -- The first part is the map area, i.e. the characters and colours.
      (X"9F20", X"00"),
      (X"9F21", X"00"),
      (X"9F22", X"10"), -- Set address to 0x00000 and increment to 1.
      (X"9F23", X"5F"), -- 0x00000
      (X"9F23", X"64"),
      (X"9F23", X"A0"),
      (X"9F23", X"64"),
      (X"9F23", X"A0"),
      (X"9F23", X"64"),
      (X"9F23", X"DF"),
      (X"9F23", X"64"),
      (X"9F23", X"20"),
      (X"9F23", X"64"),
      (X"9F23", X"20"),
      (X"9F23", X"64"),
      (X"9F23", X"20"),
      (X"9F23", X"64"),
      (X"9F23", X"E9"),
      (X"9F23", X"64"),
      (X"9F23", X"A0"), -- 0x00010
      (X"9F23", X"64"),
      (X"9F23", X"A0"),
      (X"9F23", X"64"),
      (X"9F23", X"69"),
      (X"9F23", X"64"),

      (X"9F20", X"00"),
      (X"9F21", X"01"), -- Set address to 0x00100
      (X"9F23", X"20"), -- 0x00100
      (X"9F23", X"6E"),
      (X"9F23", X"5F"),
      (X"9F23", X"6E"),
      (X"9F23", X"A0"),
      (X"9F23", X"6E"),
      (X"9F23", X"A0"),
      (X"9F23", X"6E"),
      (X"9F23", X"DF"),
      (X"9F23", X"6E"),
      (X"9F23", X"20"),
      (X"9F23", X"6E"),
      (X"9F23", X"E9"),
      (X"9F23", X"6E"),
      (X"9F23", X"A0"),
      (X"9F23", X"6E"),
      (X"9F23", X"A0"), -- 0x00110
      (X"9F23", X"6E"),
      (X"9F23", X"69"),
      (X"9F23", X"6E"),
      (X"9F23", X"20"),
      (X"9F23", X"61"),
      (X"9F23", X"20"),
      (X"9F23", X"61"),
      (X"9F23", X"2A"),
      (X"9F23", X"61"),
      (X"9F23", X"2A"),
      (X"9F23", X"61"),
      (X"9F23", X"2A"),
      (X"9F23", X"61"),
      (X"9F23", X"2A"),
      (X"9F23", X"61"),
      (X"9F23", X"20"), -- 0x00120
      (X"9F23", X"61"),
      (X"9F23", X"03"),
      (X"9F23", X"61"),
      (X"9F23", X"0F"),
      (X"9F23", X"61"),
      (X"9F23", X"0D"),
      (X"9F23", X"61"),
      (X"9F23", X"0D"),
      (X"9F23", X"61"),
      (X"9F23", X"01"),
      (X"9F23", X"61"),
      (X"9F23", X"0E"),
      (X"9F23", X"61"),
      (X"9F23", X"04"),
      (X"9F23", X"61"),
      (X"9F23", X"05"), -- 0x00130
      (X"9F23", X"61"),
      (X"9F23", X"12"),
      (X"9F23", X"61"),
      (X"9F23", X"20"),
      (X"9F23", X"61"),
      (X"9F23", X"18"),
      (X"9F23", X"61"),
      (X"9F23", X"31"),
      (X"9F23", X"61"),
      (X"9F23", X"36"),
      (X"9F23", X"61"),
      (X"9F23", X"20"),
      (X"9F23", X"61"),
      (X"9F23", X"02"),
      (X"9F23", X"61"),
      (X"9F23", X"01"), -- 0x00140
      (X"9F23", X"61"),
      (X"9F23", X"13"),
      (X"9F23", X"61"),
      (X"9F23", X"09"),
      (X"9F23", X"61"),
      (X"9F23", X"03"),
      (X"9F23", X"61"),
      (X"9F23", X"20"),
      (X"9F23", X"61"),
      (X"9F23", X"16"),
      (X"9F23", X"61"),
      (X"9F23", X"32"),
      (X"9F23", X"61"),
      (X"9F23", X"20"),
      (X"9F23", X"61"),
      (X"9F23", X"2A"), -- 0x00150
      (X"9F23", X"61"),
      (X"9F23", X"2A"),
      (X"9F23", X"61"),
      (X"9F23", X"2A"),
      (X"9F23", X"61"),
      (X"9F23", X"2A"),
      (X"9F23", X"61"),

      (X"9F20", X"00"),
      (X"9F21", X"02"), -- Set address to 0x00200
      (X"9F23", X"20"), -- 0x00200
      (X"9F23", X"63"),
      (X"9F23", X"20"),
      (X"9F23", X"63"),
      (X"9F23", X"5F"),
      (X"9F23", X"63"),
      (X"9F23", X"A0"),
      (X"9F23", X"63"),
      (X"9F23", X"A0"),
      (X"9F23", X"63"),
      (X"9F23", X"20"),
      (X"9F23", X"63"),
      (X"9F23", X"A0"),
      (X"9F23", X"63"),
      (X"9F23", X"A0"),
      (X"9F23", X"63"),
      (X"9F23", X"69"), -- 0x00210
      (X"9F23", X"63"),

      (X"9F20", X"00"),
      (X"9F21", X"03"), -- Set address to 0x00300
      (X"9F23", X"20"), -- 0x00300
      (X"9F23", X"65"),
      (X"9F23", X"20"),
      (X"9F23", X"65"),
      (X"9F23", X"20"),
      (X"9F23", X"65"),
      (X"9F23", X"20"),
      (X"9F23", X"65"),
      (X"9F23", X"A0"),
      (X"9F23", X"65"),
      (X"9F23", X"20"),
      (X"9F23", X"65"),
      (X"9F23", X"A0"),
      (X"9F23", X"65"),
      (X"9F23", X"20"),
      (X"9F23", X"61"),
      (X"9F23", X"20"), -- 0x00310
      (X"9F23", X"61"),
      (X"9F23", X"20"),
      (X"9F23", X"61"),
      (X"9F23", X"20"),
      (X"9F23", X"61"),
      (X"9F23", X"20"),
      (X"9F23", X"61"),
      (X"9F23", X"35"),
      (X"9F23", X"61"),
      (X"9F23", X"31"),
      (X"9F23", X"61"),
      (X"9F23", X"32"),
      (X"9F23", X"61"),
      (X"9F23", X"0B"),
      (X"9F23", X"61"),
      (X"9F23", X"20"), -- 0x00320
      (X"9F23", X"61"),
      (X"9F23", X"08"),
      (X"9F23", X"61"),
      (X"9F23", X"09"),
      (X"9F23", X"61"),
      (X"9F23", X"07"),
      (X"9F23", X"61"),
      (X"9F23", X"08"),
      (X"9F23", X"61"),
      (X"9F23", X"20"),
      (X"9F23", X"61"),
      (X"9F23", X"12"),
      (X"9F23", X"61"),
      (X"9F23", X"01"),
      (X"9F23", X"61"),
      (X"9F23", X"0D"), -- 0x00330
      (X"9F23", X"61"),

      (X"9F20", X"00"),
      (X"9F21", X"04"), -- Set address to 0x00400
      (X"9F23", X"20"), -- 0x00400
      (X"9F23", X"67"),
      (X"9F23", X"20"),
      (X"9F23", X"67"),
      (X"9F23", X"E9"),
      (X"9F23", X"67"),
      (X"9F23", X"A0"),
      (X"9F23", X"67"),
      (X"9F23", X"A0"),
      (X"9F23", X"67"),
      (X"9F23", X"20"),
      (X"9F23", X"67"),
      (X"9F23", X"A0"),
      (X"9F23", X"67"),
      (X"9F23", X"A0"),
      (X"9F23", X"67"),
      (X"9F23", X"DF"), -- 0x00410
      (X"9F23", X"67"),

      (X"9F20", X"00"),
      (X"9F21", X"05"), -- Set address to 0x00500
      (X"9F23", X"20"), -- 0x00500
      (X"9F23", X"68"),
      (X"9F23", X"E9"),
      (X"9F23", X"68"),
      (X"9F23", X"A0"),
      (X"9F23", X"68"),
      (X"9F23", X"A0"),
      (X"9F23", X"68"),
      (X"9F23", X"69"),
      (X"9F23", X"68"),
      (X"9F23", X"20"),
      (X"9F23", X"68"),
      (X"9F23", X"5F"),
      (X"9F23", X"68"),
      (X"9F23", X"A0"),
      (X"9F23", X"68"),
      (X"9F23", X"A0"), -- 0x00510
      (X"9F23", X"68"),
      (X"9F23", X"DF"),
      (X"9F23", X"68"),
      (X"9F23", X"20"),
      (X"9F23", X"61"),
      (X"9F23", X"20"),
      (X"9F23", X"61"),
      (X"9F23", X"33"),
      (X"9F23", X"61"),
      (X"9F23", X"38"),
      (X"9F23", X"61"),
      (X"9F23", X"36"),
      (X"9F23", X"61"),
      (X"9F23", X"35"),
      (X"9F23", X"61"),
      (X"9F23", X"35"), -- 0x00520
      (X"9F23", X"61"),
      (X"9F23", X"20"),
      (X"9F23", X"61"),
      (X"9F23", X"02"),
      (X"9F23", X"61"),
      (X"9F23", X"01"),
      (X"9F23", X"61"),
      (X"9F23", X"13"),
      (X"9F23", X"61"),
      (X"9F23", X"09"),
      (X"9F23", X"61"),
      (X"9F23", X"03"),
      (X"9F23", X"61"),
      (X"9F23", X"20"),
      (X"9F23", X"61"),
      (X"9F23", X"02"), -- 0x00530
      (X"9F23", X"61"),
      (X"9F23", X"19"),
      (X"9F23", X"61"),
      (X"9F23", X"14"),
      (X"9F23", X"61"),
      (X"9F23", X"05"),
      (X"9F23", X"61"),
      (X"9F23", X"13"),
      (X"9F23", X"61"),
      (X"9F23", X"20"),
      (X"9F23", X"61"),
      (X"9F23", X"06"),
      (X"9F23", X"61"),
      (X"9F23", X"12"),
      (X"9F23", X"61"),
      (X"9F23", X"05"), -- 0x00540
      (X"9F23", X"61"),
      (X"9F23", X"05"),
      (X"9F23", X"61"),

      (X"9F20", X"00"),
      (X"9F21", X"06"), -- Set address to 0x00600
      (X"9F23", X"E9"), -- 0x00600
      (X"9F23", X"62"),
      (X"9F23", X"A0"),
      (X"9F23", X"62"),
      (X"9F23", X"A0"),
      (X"9F23", X"62"),
      (X"9F23", X"69"),
      (X"9F23", X"62"),
      (X"9F23", X"20"),
      (X"9F23", X"62"),
      (X"9F23", X"20"),
      (X"9F23", X"62"),
      (X"9F23", X"20"),
      (X"9F23", X"62"),
      (X"9F23", X"5F"),
      (X"9F23", X"62"),
      (X"9F23", X"A0"), -- 0x00610
      (X"9F23", X"62"),
      (X"9F23", X"A0"),
      (X"9F23", X"62"),
      (X"9F23", X"DF"),
      (X"9F23", X"62"),

      (X"9F20", X"00"),
      (X"9F21", X"08"), -- Set address to 0x00800
      (X"9F23", X"12"), -- 0x00800
      (X"9F23", X"61"),
      (X"9F23", X"05"),
      (X"9F23", X"61"),
      (X"9F23", X"01"),
      (X"9F23", X"61"),
      (X"9F23", X"04"),
      (X"9F23", X"61"),
      (X"9F23", X"19"),
      (X"9F23", X"61"),
      (X"9F23", X"2E"),
      (X"9F23", X"61"),

      -- The second part is the tile map, i.e. the font
      (X"9F20", X"00"),
      (X"9F21", X"F8"), -- Set address to 0x0F800
      (X"9F23", X"3C"), -- 0x0F800
      (X"9F23", X"66"),
      (X"9F23", X"6E"),
      (X"9F23", X"6E"),
      (X"9F23", X"60"),
      (X"9F23", X"62"),
      (X"9F23", X"3C"),
      (X"9F23", X"00"),
      (X"9F23", X"18"),
      (X"9F23", X"3C"),
      (X"9F23", X"66"),
      (X"9F23", X"7E"),
      (X"9F23", X"66"),
      (X"9F23", X"66"),
      (X"9F23", X"66"),
      (X"9F23", X"00"),
      (X"9F23", X"7C"),
      (X"9F23", X"66"),
      (X"9F23", X"66"),
      (X"9F23", X"7C"),
      (X"9F23", X"66"),
      (X"9F23", X"66"),
      (X"9F23", X"7C"),
      (X"9F23", X"00"),
      (X"9F23", X"3C"),
      (X"9F23", X"66"),
      (X"9F23", X"60"),
      (X"9F23", X"60"),
      (X"9F23", X"60"),
      (X"9F23", X"66"),
      (X"9F23", X"3C"),
      (X"9F23", X"00"),
      (X"9F23", X"78"),
      (X"9F23", X"6C"),
      (X"9F23", X"66"),
      (X"9F23", X"66"),
      (X"9F23", X"66"),
      (X"9F23", X"6C"),
      (X"9F23", X"78"),
      (X"9F23", X"00"),
      (X"9F23", X"7E"),
      (X"9F23", X"60"),
      (X"9F23", X"60"),
      (X"9F23", X"78"),
      (X"9F23", X"60"),
      (X"9F23", X"60"),
      (X"9F23", X"7E"),
      (X"9F23", X"00"),
      (X"9F23", X"7E"),
      (X"9F23", X"60"),
      (X"9F23", X"60"),
      (X"9F23", X"78"),
      (X"9F23", X"60"),
      (X"9F23", X"60"),
      (X"9F23", X"60"),
      (X"9F23", X"00"),
      (X"9F23", X"3C"),
      (X"9F23", X"66"),
      (X"9F23", X"60"),
      (X"9F23", X"6E"),
      (X"9F23", X"66"),
      (X"9F23", X"66"),
      (X"9F23", X"3C"),
      (X"9F23", X"00"),
      (X"9F23", X"66"),
      (X"9F23", X"66"),
      (X"9F23", X"66"),
      (X"9F23", X"7E"),
      (X"9F23", X"66"),
      (X"9F23", X"66"),
      (X"9F23", X"66"),
      (X"9F23", X"00"),
      (X"9F23", X"3C"),
      (X"9F23", X"18"),
      (X"9F23", X"18"),
      (X"9F23", X"18"),
      (X"9F23", X"18"),
      (X"9F23", X"18"),
      (X"9F23", X"3C"),
      (X"9F23", X"00"),
      (X"9F23", X"1E"),
      (X"9F23", X"0C"),
      (X"9F23", X"0C"),
      (X"9F23", X"0C"),
      (X"9F23", X"0C"),
      (X"9F23", X"6C"),
      (X"9F23", X"38"),
      (X"9F23", X"00"),
      (X"9F23", X"66"),
      (X"9F23", X"6C"),
      (X"9F23", X"78"),
      (X"9F23", X"70"),
      (X"9F23", X"78"),
      (X"9F23", X"6C"),
      (X"9F23", X"66"),
      (X"9F23", X"00"),
      (X"9F23", X"60"),
      (X"9F23", X"60"),
      (X"9F23", X"60"),
      (X"9F23", X"60"),
      (X"9F23", X"60"),
      (X"9F23", X"60"),
      (X"9F23", X"7E"),
      (X"9F23", X"00"),
      (X"9F23", X"63"),
      (X"9F23", X"77"),
      (X"9F23", X"7F"),
      (X"9F23", X"6B"),
      (X"9F23", X"63"),
      (X"9F23", X"63"),
      (X"9F23", X"63"),
      (X"9F23", X"00"),
      (X"9F23", X"66"),
      (X"9F23", X"76"),
      (X"9F23", X"7E"),
      (X"9F23", X"7E"),
      (X"9F23", X"6E"),
      (X"9F23", X"66"),
      (X"9F23", X"66"),
      (X"9F23", X"00"),
      (X"9F23", X"3C"),
      (X"9F23", X"66"),
      (X"9F23", X"66"),
      (X"9F23", X"66"),
      (X"9F23", X"66"),
      (X"9F23", X"66"),
      (X"9F23", X"3C"),
      (X"9F23", X"00"),
      (X"9F23", X"7C"),
      (X"9F23", X"66"),
      (X"9F23", X"66"),
      (X"9F23", X"7C"),
      (X"9F23", X"60"),
      (X"9F23", X"60"),
      (X"9F23", X"60"),
      (X"9F23", X"00"),
      (X"9F23", X"3C"),
      (X"9F23", X"66"),
      (X"9F23", X"66"),
      (X"9F23", X"66"),
      (X"9F23", X"66"),
      (X"9F23", X"3C"),
      (X"9F23", X"0E"),
      (X"9F23", X"00"),
      (X"9F23", X"7C"),
      (X"9F23", X"66"),
      (X"9F23", X"66"),
      (X"9F23", X"7C"),
      (X"9F23", X"78"),
      (X"9F23", X"6C"),
      (X"9F23", X"66"),
      (X"9F23", X"00"),
      (X"9F23", X"3C"),
      (X"9F23", X"66"),
      (X"9F23", X"60"),
      (X"9F23", X"3C"),
      (X"9F23", X"06"),
      (X"9F23", X"66"),
      (X"9F23", X"3C"),
      (X"9F23", X"00"),
      (X"9F23", X"7E"),
      (X"9F23", X"18"),
      (X"9F23", X"18"),
      (X"9F23", X"18"),
      (X"9F23", X"18"),
      (X"9F23", X"18"),
      (X"9F23", X"18"),
      (X"9F23", X"00"),
      (X"9F23", X"66"),
      (X"9F23", X"66"),
      (X"9F23", X"66"),
      (X"9F23", X"66"),
      (X"9F23", X"66"),
      (X"9F23", X"66"),
      (X"9F23", X"3C"),
      (X"9F23", X"00"),
      (X"9F23", X"66"),
      (X"9F23", X"66"),
      (X"9F23", X"66"),
      (X"9F23", X"66"),
      (X"9F23", X"66"),
      (X"9F23", X"3C"),
      (X"9F23", X"18"),
      (X"9F23", X"00"),
      (X"9F23", X"63"),
      (X"9F23", X"63"),
      (X"9F23", X"63"),
      (X"9F23", X"6B"),
      (X"9F23", X"7F"),
      (X"9F23", X"77"),
      (X"9F23", X"63"),
      (X"9F23", X"00"),
      (X"9F23", X"66"),
      (X"9F23", X"66"),
      (X"9F23", X"3C"),
      (X"9F23", X"18"),
      (X"9F23", X"3C"),
      (X"9F23", X"66"),
      (X"9F23", X"66"),
      (X"9F23", X"00"),
      (X"9F23", X"66"),
      (X"9F23", X"66"),
      (X"9F23", X"66"),
      (X"9F23", X"3C"),
      (X"9F23", X"18"),
      (X"9F23", X"18"),
      (X"9F23", X"18"),
      (X"9F23", X"00"),
      (X"9F23", X"7E"),
      (X"9F23", X"06"),
      (X"9F23", X"0C"),
      (X"9F23", X"18"),
      (X"9F23", X"30"),
      (X"9F23", X"60"),
      (X"9F23", X"7E"),
      (X"9F23", X"00"),
      (X"9F23", X"3C"),
      (X"9F23", X"30"),
      (X"9F23", X"30"),
      (X"9F23", X"30"),
      (X"9F23", X"30"),
      (X"9F23", X"30"),
      (X"9F23", X"3C"),
      (X"9F23", X"00"),
      (X"9F23", X"0C"),
      (X"9F23", X"12"),
      (X"9F23", X"30"),
      (X"9F23", X"7C"),
      (X"9F23", X"30"),
      (X"9F23", X"62"),
      (X"9F23", X"FC"),
      (X"9F23", X"00"),
      (X"9F23", X"3C"),
      (X"9F23", X"0C"),
      (X"9F23", X"0C"),
      (X"9F23", X"0C"),
      (X"9F23", X"0C"),
      (X"9F23", X"0C"),
      (X"9F23", X"3C"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"18"),
      (X"9F23", X"3C"),
      (X"9F23", X"7E"),
      (X"9F23", X"18"),
      (X"9F23", X"18"),
      (X"9F23", X"18"),
      (X"9F23", X"18"),
      (X"9F23", X"00"),
      (X"9F23", X"10"),
      (X"9F23", X"30"),
      (X"9F23", X"7F"),
      (X"9F23", X"7F"),
      (X"9F23", X"30"),
      (X"9F23", X"10"),
      (X"9F23", X"00"),
      (X"9F23", X"00"), -- 0x0F900
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"18"),
      (X"9F23", X"18"),
      (X"9F23", X"18"),
      (X"9F23", X"18"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"18"),
      (X"9F23", X"00"),
      (X"9F23", X"66"),
      (X"9F23", X"66"),
      (X"9F23", X"66"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"66"),
      (X"9F23", X"66"),
      (X"9F23", X"FF"),
      (X"9F23", X"66"),
      (X"9F23", X"FF"),
      (X"9F23", X"66"),
      (X"9F23", X"66"),
      (X"9F23", X"00"),
      (X"9F23", X"18"),
      (X"9F23", X"3E"),
      (X"9F23", X"60"),
      (X"9F23", X"3C"),
      (X"9F23", X"06"),
      (X"9F23", X"7C"),
      (X"9F23", X"18"),
      (X"9F23", X"00"),
      (X"9F23", X"62"),
      (X"9F23", X"66"),
      (X"9F23", X"0C"),
      (X"9F23", X"18"),
      (X"9F23", X"30"),
      (X"9F23", X"66"),
      (X"9F23", X"46"),
      (X"9F23", X"00"),
      (X"9F23", X"3C"),
      (X"9F23", X"66"),
      (X"9F23", X"3C"),
      (X"9F23", X"38"),
      (X"9F23", X"67"),
      (X"9F23", X"66"),
      (X"9F23", X"3F"),
      (X"9F23", X"00"),
      (X"9F23", X"06"),
      (X"9F23", X"0C"),
      (X"9F23", X"18"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"0C"),
      (X"9F23", X"18"),
      (X"9F23", X"30"),
      (X"9F23", X"30"),
      (X"9F23", X"30"),
      (X"9F23", X"18"),
      (X"9F23", X"0C"),
      (X"9F23", X"00"),
      (X"9F23", X"30"),
      (X"9F23", X"18"),
      (X"9F23", X"0C"),
      (X"9F23", X"0C"),
      (X"9F23", X"0C"),
      (X"9F23", X"18"),
      (X"9F23", X"30"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"66"),
      (X"9F23", X"3C"),
      (X"9F23", X"FF"),
      (X"9F23", X"3C"),
      (X"9F23", X"66"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"18"),
      (X"9F23", X"18"),
      (X"9F23", X"7E"),
      (X"9F23", X"18"),
      (X"9F23", X"18"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"18"),
      (X"9F23", X"18"),
      (X"9F23", X"30"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"7E"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"18"),
      (X"9F23", X"18"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"03"),
      (X"9F23", X"06"),
      (X"9F23", X"0C"),
      (X"9F23", X"18"),
      (X"9F23", X"30"),
      (X"9F23", X"60"),
      (X"9F23", X"00"),
      (X"9F23", X"3C"),
      (X"9F23", X"66"),
      (X"9F23", X"6E"),
      (X"9F23", X"76"),
      (X"9F23", X"66"),
      (X"9F23", X"66"),
      (X"9F23", X"3C"),
      (X"9F23", X"00"),
      (X"9F23", X"18"),
      (X"9F23", X"18"),
      (X"9F23", X"38"),
      (X"9F23", X"18"),
      (X"9F23", X"18"),
      (X"9F23", X"18"),
      (X"9F23", X"7E"),
      (X"9F23", X"00"),
      (X"9F23", X"3C"),
      (X"9F23", X"66"),
      (X"9F23", X"06"),
      (X"9F23", X"0C"),
      (X"9F23", X"30"),
      (X"9F23", X"60"),
      (X"9F23", X"7E"),
      (X"9F23", X"00"),
      (X"9F23", X"3C"),
      (X"9F23", X"66"),
      (X"9F23", X"06"),
      (X"9F23", X"1C"),
      (X"9F23", X"06"),
      (X"9F23", X"66"),
      (X"9F23", X"3C"),
      (X"9F23", X"00"),
      (X"9F23", X"06"),
      (X"9F23", X"0E"),
      (X"9F23", X"1E"),
      (X"9F23", X"66"),
      (X"9F23", X"7F"),
      (X"9F23", X"06"),
      (X"9F23", X"06"),
      (X"9F23", X"00"),
      (X"9F23", X"7E"),
      (X"9F23", X"60"),
      (X"9F23", X"7C"),
      (X"9F23", X"06"),
      (X"9F23", X"06"),
      (X"9F23", X"66"),
      (X"9F23", X"3C"),
      (X"9F23", X"00"),
      (X"9F23", X"3C"),
      (X"9F23", X"66"),
      (X"9F23", X"60"),
      (X"9F23", X"7C"),
      (X"9F23", X"66"),
      (X"9F23", X"66"),
      (X"9F23", X"3C"),
      (X"9F23", X"00"),
      (X"9F23", X"7E"),
      (X"9F23", X"66"),
      (X"9F23", X"0C"),
      (X"9F23", X"18"),
      (X"9F23", X"18"),
      (X"9F23", X"18"),
      (X"9F23", X"18"),
      (X"9F23", X"00"),
      (X"9F23", X"3C"),
      (X"9F23", X"66"),
      (X"9F23", X"66"),
      (X"9F23", X"3C"),
      (X"9F23", X"66"),
      (X"9F23", X"66"),
      (X"9F23", X"3C"),
      (X"9F23", X"00"),
      (X"9F23", X"3C"),
      (X"9F23", X"66"),
      (X"9F23", X"66"),
      (X"9F23", X"3E"),
      (X"9F23", X"06"),
      (X"9F23", X"66"),
      (X"9F23", X"3C"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"18"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"18"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"18"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"18"),
      (X"9F23", X"18"),
      (X"9F23", X"30"),
      (X"9F23", X"0E"),
      (X"9F23", X"18"),
      (X"9F23", X"30"),
      (X"9F23", X"60"),
      (X"9F23", X"30"),
      (X"9F23", X"18"),
      (X"9F23", X"0E"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"7E"),
      (X"9F23", X"00"),
      (X"9F23", X"7E"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"70"),
      (X"9F23", X"18"),
      (X"9F23", X"0C"),
      (X"9F23", X"06"),
      (X"9F23", X"0C"),
      (X"9F23", X"18"),
      (X"9F23", X"70"),
      (X"9F23", X"00"),
      (X"9F23", X"3C"),
      (X"9F23", X"66"),
      (X"9F23", X"06"),
      (X"9F23", X"0C"),
      (X"9F23", X"18"),
      (X"9F23", X"00"),
      (X"9F23", X"18"),
      (X"9F23", X"00"),
      (X"9F23", X"00"), -- 0x0FA00
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"08"),
      (X"9F23", X"1C"),
      (X"9F23", X"3E"),
      (X"9F23", X"7F"),
      (X"9F23", X"7F"),
      (X"9F23", X"1C"),
      (X"9F23", X"3E"),
      (X"9F23", X"00"),
      (X"9F23", X"18"),
      (X"9F23", X"18"),
      (X"9F23", X"18"),
      (X"9F23", X"18"),
      (X"9F23", X"18"),
      (X"9F23", X"18"),
      (X"9F23", X"18"),
      (X"9F23", X"18"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"30"),
      (X"9F23", X"30"),
      (X"9F23", X"30"),
      (X"9F23", X"30"),
      (X"9F23", X"30"),
      (X"9F23", X"30"),
      (X"9F23", X"30"),
      (X"9F23", X"30"),
      (X"9F23", X"0C"),
      (X"9F23", X"0C"),
      (X"9F23", X"0C"),
      (X"9F23", X"0C"),
      (X"9F23", X"0C"),
      (X"9F23", X"0C"),
      (X"9F23", X"0C"),
      (X"9F23", X"0C"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"E0"),
      (X"9F23", X"F0"),
      (X"9F23", X"38"),
      (X"9F23", X"18"),
      (X"9F23", X"18"),
      (X"9F23", X"18"),
      (X"9F23", X"18"),
      (X"9F23", X"1C"),
      (X"9F23", X"0F"),
      (X"9F23", X"07"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"18"),
      (X"9F23", X"18"),
      (X"9F23", X"38"),
      (X"9F23", X"F0"),
      (X"9F23", X"E0"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"C0"),
      (X"9F23", X"C0"),
      (X"9F23", X"C0"),
      (X"9F23", X"C0"),
      (X"9F23", X"C0"),
      (X"9F23", X"C0"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"C0"),
      (X"9F23", X"E0"),
      (X"9F23", X"70"),
      (X"9F23", X"38"),
      (X"9F23", X"1C"),
      (X"9F23", X"0E"),
      (X"9F23", X"07"),
      (X"9F23", X"03"),
      (X"9F23", X"03"),
      (X"9F23", X"07"),
      (X"9F23", X"0E"),
      (X"9F23", X"1C"),
      (X"9F23", X"38"),
      (X"9F23", X"70"),
      (X"9F23", X"E0"),
      (X"9F23", X"C0"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"C0"),
      (X"9F23", X"C0"),
      (X"9F23", X"C0"),
      (X"9F23", X"C0"),
      (X"9F23", X"C0"),
      (X"9F23", X"C0"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"03"),
      (X"9F23", X"03"),
      (X"9F23", X"03"),
      (X"9F23", X"03"),
      (X"9F23", X"03"),
      (X"9F23", X"03"),
      (X"9F23", X"00"),
      (X"9F23", X"3C"),
      (X"9F23", X"7E"),
      (X"9F23", X"7E"),
      (X"9F23", X"7E"),
      (X"9F23", X"7E"),
      (X"9F23", X"3C"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"00"),
      (X"9F23", X"36"),
      (X"9F23", X"7F"),
      (X"9F23", X"7F"),
      (X"9F23", X"7F"),
      (X"9F23", X"3E"),
      (X"9F23", X"1C"),
      (X"9F23", X"08"),
      (X"9F23", X"00"),
      (X"9F23", X"60"),
      (X"9F23", X"60"),
      (X"9F23", X"60"),
      (X"9F23", X"60"),
      (X"9F23", X"60"),
      (X"9F23", X"60"),
      (X"9F23", X"60"),
      (X"9F23", X"60"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"07"),
      (X"9F23", X"0F"),
      (X"9F23", X"1C"),
      (X"9F23", X"18"),
      (X"9F23", X"18"),
      (X"9F23", X"C3"),
      (X"9F23", X"E7"),
      (X"9F23", X"7E"),
      (X"9F23", X"3C"),
      (X"9F23", X"3C"),
      (X"9F23", X"7E"),
      (X"9F23", X"E7"),
      (X"9F23", X"C3"),
      (X"9F23", X"00"),
      (X"9F23", X"3C"),
      (X"9F23", X"7E"),
      (X"9F23", X"66"),
      (X"9F23", X"66"),
      (X"9F23", X"7E"),
      (X"9F23", X"3C"),
      (X"9F23", X"00"),
      (X"9F23", X"18"),
      (X"9F23", X"18"),
      (X"9F23", X"66"),
      (X"9F23", X"66"),
      (X"9F23", X"18"),
      (X"9F23", X"18"),
      (X"9F23", X"3C"),
      (X"9F23", X"00"),
      (X"9F23", X"06"),
      (X"9F23", X"06"),
      (X"9F23", X"06"),
      (X"9F23", X"06"),
      (X"9F23", X"06"),
      (X"9F23", X"06"),
      (X"9F23", X"06"),
      (X"9F23", X"06"),
      (X"9F23", X"08"),
      (X"9F23", X"1C"),
      (X"9F23", X"3E"),
      (X"9F23", X"7F"),
      (X"9F23", X"3E"),
      (X"9F23", X"1C"),
      (X"9F23", X"08"),
      (X"9F23", X"00"),
      (X"9F23", X"18"),
      (X"9F23", X"18"),
      (X"9F23", X"18"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"18"),
      (X"9F23", X"18"),
      (X"9F23", X"18"),
      (X"9F23", X"C0"),
      (X"9F23", X"C0"),
      (X"9F23", X"30"),
      (X"9F23", X"30"),
      (X"9F23", X"C0"),
      (X"9F23", X"C0"),
      (X"9F23", X"30"),
      (X"9F23", X"30"),
      (X"9F23", X"18"),
      (X"9F23", X"18"),
      (X"9F23", X"18"),
      (X"9F23", X"18"),
      (X"9F23", X"18"),
      (X"9F23", X"18"),
      (X"9F23", X"18"),
      (X"9F23", X"18"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"03"),
      (X"9F23", X"3E"),
      (X"9F23", X"76"),
      (X"9F23", X"36"),
      (X"9F23", X"36"),
      (X"9F23", X"00"),
      (X"9F23", X"FF"),
      (X"9F23", X"7F"),
      (X"9F23", X"3F"),
      (X"9F23", X"1F"),
      (X"9F23", X"0F"),
      (X"9F23", X"07"),
      (X"9F23", X"03"),
      (X"9F23", X"01"),
      (X"9F23", X"00"), -- 0x0FB00
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"F0"),
      (X"9F23", X"F0"),
      (X"9F23", X"F0"),
      (X"9F23", X"F0"),
      (X"9F23", X"F0"),
      (X"9F23", X"F0"),
      (X"9F23", X"F0"),
      (X"9F23", X"F0"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"FF"),
      (X"9F23", X"C0"),
      (X"9F23", X"C0"),
      (X"9F23", X"C0"),
      (X"9F23", X"C0"),
      (X"9F23", X"C0"),
      (X"9F23", X"C0"),
      (X"9F23", X"C0"),
      (X"9F23", X"C0"),
      (X"9F23", X"CC"),
      (X"9F23", X"CC"),
      (X"9F23", X"33"),
      (X"9F23", X"33"),
      (X"9F23", X"CC"),
      (X"9F23", X"CC"),
      (X"9F23", X"33"),
      (X"9F23", X"33"),
      (X"9F23", X"03"),
      (X"9F23", X"03"),
      (X"9F23", X"03"),
      (X"9F23", X"03"),
      (X"9F23", X"03"),
      (X"9F23", X"03"),
      (X"9F23", X"03"),
      (X"9F23", X"03"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"CC"),
      (X"9F23", X"CC"),
      (X"9F23", X"33"),
      (X"9F23", X"33"),
      (X"9F23", X"FF"),
      (X"9F23", X"FE"),
      (X"9F23", X"FC"),
      (X"9F23", X"F8"),
      (X"9F23", X"F0"),
      (X"9F23", X"E0"),
      (X"9F23", X"C0"),
      (X"9F23", X"80"),
      (X"9F23", X"03"),
      (X"9F23", X"03"),
      (X"9F23", X"03"),
      (X"9F23", X"03"),
      (X"9F23", X"03"),
      (X"9F23", X"03"),
      (X"9F23", X"03"),
      (X"9F23", X"03"),
      (X"9F23", X"18"),
      (X"9F23", X"18"),
      (X"9F23", X"18"),
      (X"9F23", X"1F"),
      (X"9F23", X"1F"),
      (X"9F23", X"18"),
      (X"9F23", X"18"),
      (X"9F23", X"18"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"0F"),
      (X"9F23", X"0F"),
      (X"9F23", X"0F"),
      (X"9F23", X"0F"),
      (X"9F23", X"18"),
      (X"9F23", X"18"),
      (X"9F23", X"18"),
      (X"9F23", X"1F"),
      (X"9F23", X"1F"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"F8"),
      (X"9F23", X"F8"),
      (X"9F23", X"18"),
      (X"9F23", X"18"),
      (X"9F23", X"18"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"1F"),
      (X"9F23", X"1F"),
      (X"9F23", X"18"),
      (X"9F23", X"18"),
      (X"9F23", X"18"),
      (X"9F23", X"18"),
      (X"9F23", X"18"),
      (X"9F23", X"18"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"18"),
      (X"9F23", X"18"),
      (X"9F23", X"18"),
      (X"9F23", X"18"),
      (X"9F23", X"18"),
      (X"9F23", X"18"),
      (X"9F23", X"F8"),
      (X"9F23", X"F8"),
      (X"9F23", X"18"),
      (X"9F23", X"18"),
      (X"9F23", X"18"),
      (X"9F23", X"C0"),
      (X"9F23", X"C0"),
      (X"9F23", X"C0"),
      (X"9F23", X"C0"),
      (X"9F23", X"C0"),
      (X"9F23", X"C0"),
      (X"9F23", X"C0"),
      (X"9F23", X"C0"),
      (X"9F23", X"E0"),
      (X"9F23", X"E0"),
      (X"9F23", X"E0"),
      (X"9F23", X"E0"),
      (X"9F23", X"E0"),
      (X"9F23", X"E0"),
      (X"9F23", X"E0"),
      (X"9F23", X"E0"),
      (X"9F23", X"07"),
      (X"9F23", X"07"),
      (X"9F23", X"07"),
      (X"9F23", X"07"),
      (X"9F23", X"07"),
      (X"9F23", X"07"),
      (X"9F23", X"07"),
      (X"9F23", X"07"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"03"),
      (X"9F23", X"03"),
      (X"9F23", X"03"),
      (X"9F23", X"03"),
      (X"9F23", X"03"),
      (X"9F23", X"03"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"F0"),
      (X"9F23", X"F0"),
      (X"9F23", X"F0"),
      (X"9F23", X"F0"),
      (X"9F23", X"0F"),
      (X"9F23", X"0F"),
      (X"9F23", X"0F"),
      (X"9F23", X"0F"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"18"),
      (X"9F23", X"18"),
      (X"9F23", X"18"),
      (X"9F23", X"F8"),
      (X"9F23", X"F8"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"F0"),
      (X"9F23", X"F0"),
      (X"9F23", X"F0"),
      (X"9F23", X"F0"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"F0"),
      (X"9F23", X"F0"),
      (X"9F23", X"F0"),
      (X"9F23", X"F0"),
      (X"9F23", X"0F"),
      (X"9F23", X"0F"),
      (X"9F23", X"0F"),
      (X"9F23", X"0F"),
      (X"9F23", X"C3"), -- 0x0FC00
      (X"9F23", X"99"),
      (X"9F23", X"91"),
      (X"9F23", X"91"),
      (X"9F23", X"9F"),
      (X"9F23", X"9D"),
      (X"9F23", X"C3"),
      (X"9F23", X"FF"),
      (X"9F23", X"E7"),
      (X"9F23", X"C3"),
      (X"9F23", X"99"),
      (X"9F23", X"81"),
      (X"9F23", X"99"),
      (X"9F23", X"99"),
      (X"9F23", X"99"),
      (X"9F23", X"FF"),
      (X"9F23", X"83"),
      (X"9F23", X"99"),
      (X"9F23", X"99"),
      (X"9F23", X"83"),
      (X"9F23", X"99"),
      (X"9F23", X"99"),
      (X"9F23", X"83"),
      (X"9F23", X"FF"),
      (X"9F23", X"C3"),
      (X"9F23", X"99"),
      (X"9F23", X"9F"),
      (X"9F23", X"9F"),
      (X"9F23", X"9F"),
      (X"9F23", X"99"),
      (X"9F23", X"C3"),
      (X"9F23", X"FF"),
      (X"9F23", X"87"),
      (X"9F23", X"93"),
      (X"9F23", X"99"),
      (X"9F23", X"99"),
      (X"9F23", X"99"),
      (X"9F23", X"93"),
      (X"9F23", X"87"),
      (X"9F23", X"FF"),
      (X"9F23", X"81"),
      (X"9F23", X"9F"),
      (X"9F23", X"9F"),
      (X"9F23", X"87"),
      (X"9F23", X"9F"),
      (X"9F23", X"9F"),
      (X"9F23", X"81"),
      (X"9F23", X"FF"),
      (X"9F23", X"81"),
      (X"9F23", X"9F"),
      (X"9F23", X"9F"),
      (X"9F23", X"87"),
      (X"9F23", X"9F"),
      (X"9F23", X"9F"),
      (X"9F23", X"9F"),
      (X"9F23", X"FF"),
      (X"9F23", X"C3"),
      (X"9F23", X"99"),
      (X"9F23", X"9F"),
      (X"9F23", X"91"),
      (X"9F23", X"99"),
      (X"9F23", X"99"),
      (X"9F23", X"C3"),
      (X"9F23", X"FF"),
      (X"9F23", X"99"),
      (X"9F23", X"99"),
      (X"9F23", X"99"),
      (X"9F23", X"81"),
      (X"9F23", X"99"),
      (X"9F23", X"99"),
      (X"9F23", X"99"),
      (X"9F23", X"FF"),
      (X"9F23", X"C3"),
      (X"9F23", X"E7"),
      (X"9F23", X"E7"),
      (X"9F23", X"E7"),
      (X"9F23", X"E7"),
      (X"9F23", X"E7"),
      (X"9F23", X"C3"),
      (X"9F23", X"FF"),
      (X"9F23", X"E1"),
      (X"9F23", X"F3"),
      (X"9F23", X"F3"),
      (X"9F23", X"F3"),
      (X"9F23", X"F3"),
      (X"9F23", X"93"),
      (X"9F23", X"C7"),
      (X"9F23", X"FF"),
      (X"9F23", X"99"),
      (X"9F23", X"93"),
      (X"9F23", X"87"),
      (X"9F23", X"8F"),
      (X"9F23", X"87"),
      (X"9F23", X"93"),
      (X"9F23", X"99"),
      (X"9F23", X"FF"),
      (X"9F23", X"9F"),
      (X"9F23", X"9F"),
      (X"9F23", X"9F"),
      (X"9F23", X"9F"),
      (X"9F23", X"9F"),
      (X"9F23", X"9F"),
      (X"9F23", X"81"),
      (X"9F23", X"FF"),
      (X"9F23", X"9C"),
      (X"9F23", X"88"),
      (X"9F23", X"80"),
      (X"9F23", X"94"),
      (X"9F23", X"9C"),
      (X"9F23", X"9C"),
      (X"9F23", X"9C"),
      (X"9F23", X"FF"),
      (X"9F23", X"99"),
      (X"9F23", X"89"),
      (X"9F23", X"81"),
      (X"9F23", X"81"),
      (X"9F23", X"91"),
      (X"9F23", X"99"),
      (X"9F23", X"99"),
      (X"9F23", X"FF"),
      (X"9F23", X"C3"),
      (X"9F23", X"99"),
      (X"9F23", X"99"),
      (X"9F23", X"99"),
      (X"9F23", X"99"),
      (X"9F23", X"99"),
      (X"9F23", X"C3"),
      (X"9F23", X"FF"),
      (X"9F23", X"83"),
      (X"9F23", X"99"),
      (X"9F23", X"99"),
      (X"9F23", X"83"),
      (X"9F23", X"9F"),
      (X"9F23", X"9F"),
      (X"9F23", X"9F"),
      (X"9F23", X"FF"),
      (X"9F23", X"C3"),
      (X"9F23", X"99"),
      (X"9F23", X"99"),
      (X"9F23", X"99"),
      (X"9F23", X"99"),
      (X"9F23", X"C3"),
      (X"9F23", X"F1"),
      (X"9F23", X"FF"),
      (X"9F23", X"83"),
      (X"9F23", X"99"),
      (X"9F23", X"99"),
      (X"9F23", X"83"),
      (X"9F23", X"87"),
      (X"9F23", X"93"),
      (X"9F23", X"99"),
      (X"9F23", X"FF"),
      (X"9F23", X"C3"),
      (X"9F23", X"99"),
      (X"9F23", X"9F"),
      (X"9F23", X"C3"),
      (X"9F23", X"F9"),
      (X"9F23", X"99"),
      (X"9F23", X"C3"),
      (X"9F23", X"FF"),
      (X"9F23", X"81"),
      (X"9F23", X"E7"),
      (X"9F23", X"E7"),
      (X"9F23", X"E7"),
      (X"9F23", X"E7"),
      (X"9F23", X"E7"),
      (X"9F23", X"E7"),
      (X"9F23", X"FF"),
      (X"9F23", X"99"),
      (X"9F23", X"99"),
      (X"9F23", X"99"),
      (X"9F23", X"99"),
      (X"9F23", X"99"),
      (X"9F23", X"99"),
      (X"9F23", X"C3"),
      (X"9F23", X"FF"),
      (X"9F23", X"99"),
      (X"9F23", X"99"),
      (X"9F23", X"99"),
      (X"9F23", X"99"),
      (X"9F23", X"99"),
      (X"9F23", X"C3"),
      (X"9F23", X"E7"),
      (X"9F23", X"FF"),
      (X"9F23", X"9C"),
      (X"9F23", X"9C"),
      (X"9F23", X"9C"),
      (X"9F23", X"94"),
      (X"9F23", X"80"),
      (X"9F23", X"88"),
      (X"9F23", X"9C"),
      (X"9F23", X"FF"),
      (X"9F23", X"99"),
      (X"9F23", X"99"),
      (X"9F23", X"C3"),
      (X"9F23", X"E7"),
      (X"9F23", X"C3"),
      (X"9F23", X"99"),
      (X"9F23", X"99"),
      (X"9F23", X"FF"),
      (X"9F23", X"99"),
      (X"9F23", X"99"),
      (X"9F23", X"99"),
      (X"9F23", X"C3"),
      (X"9F23", X"E7"),
      (X"9F23", X"E7"),
      (X"9F23", X"E7"),
      (X"9F23", X"FF"),
      (X"9F23", X"81"),
      (X"9F23", X"F9"),
      (X"9F23", X"F3"),
      (X"9F23", X"E7"),
      (X"9F23", X"CF"),
      (X"9F23", X"9F"),
      (X"9F23", X"81"),
      (X"9F23", X"FF"),
      (X"9F23", X"C3"),
      (X"9F23", X"CF"),
      (X"9F23", X"CF"),
      (X"9F23", X"CF"),
      (X"9F23", X"CF"),
      (X"9F23", X"CF"),
      (X"9F23", X"C3"),
      (X"9F23", X"FF"),
      (X"9F23", X"F3"),
      (X"9F23", X"ED"),
      (X"9F23", X"CF"),
      (X"9F23", X"83"),
      (X"9F23", X"CF"),
      (X"9F23", X"9D"),
      (X"9F23", X"03"),
      (X"9F23", X"FF"),
      (X"9F23", X"C3"),
      (X"9F23", X"F3"),
      (X"9F23", X"F3"),
      (X"9F23", X"F3"),
      (X"9F23", X"F3"),
      (X"9F23", X"F3"),
      (X"9F23", X"C3"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"E7"),
      (X"9F23", X"C3"),
      (X"9F23", X"81"),
      (X"9F23", X"E7"),
      (X"9F23", X"E7"),
      (X"9F23", X"E7"),
      (X"9F23", X"E7"),
      (X"9F23", X"FF"),
      (X"9F23", X"EF"),
      (X"9F23", X"CF"),
      (X"9F23", X"80"),
      (X"9F23", X"80"),
      (X"9F23", X"CF"),
      (X"9F23", X"EF"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"), -- 0x0FD00
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"E7"),
      (X"9F23", X"E7"),
      (X"9F23", X"E7"),
      (X"9F23", X"E7"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"E7"),
      (X"9F23", X"FF"),
      (X"9F23", X"99"),
      (X"9F23", X"99"),
      (X"9F23", X"99"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"99"),
      (X"9F23", X"99"),
      (X"9F23", X"00"),
      (X"9F23", X"99"),
      (X"9F23", X"00"),
      (X"9F23", X"99"),
      (X"9F23", X"99"),
      (X"9F23", X"FF"),
      (X"9F23", X"E7"),
      (X"9F23", X"C1"),
      (X"9F23", X"9F"),
      (X"9F23", X"C3"),
      (X"9F23", X"F9"),
      (X"9F23", X"83"),
      (X"9F23", X"E7"),
      (X"9F23", X"FF"),
      (X"9F23", X"9D"),
      (X"9F23", X"99"),
      (X"9F23", X"F3"),
      (X"9F23", X"E7"),
      (X"9F23", X"CF"),
      (X"9F23", X"99"),
      (X"9F23", X"B9"),
      (X"9F23", X"FF"),
      (X"9F23", X"C3"),
      (X"9F23", X"99"),
      (X"9F23", X"C3"),
      (X"9F23", X"C7"),
      (X"9F23", X"98"),
      (X"9F23", X"99"),
      (X"9F23", X"C0"),
      (X"9F23", X"FF"),
      (X"9F23", X"F9"),
      (X"9F23", X"F3"),
      (X"9F23", X"E7"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"F3"),
      (X"9F23", X"E7"),
      (X"9F23", X"CF"),
      (X"9F23", X"CF"),
      (X"9F23", X"CF"),
      (X"9F23", X"E7"),
      (X"9F23", X"F3"),
      (X"9F23", X"FF"),
      (X"9F23", X"CF"),
      (X"9F23", X"E7"),
      (X"9F23", X"F3"),
      (X"9F23", X"F3"),
      (X"9F23", X"F3"),
      (X"9F23", X"E7"),
      (X"9F23", X"CF"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"99"),
      (X"9F23", X"C3"),
      (X"9F23", X"00"),
      (X"9F23", X"C3"),
      (X"9F23", X"99"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"E7"),
      (X"9F23", X"E7"),
      (X"9F23", X"81"),
      (X"9F23", X"E7"),
      (X"9F23", X"E7"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"E7"),
      (X"9F23", X"E7"),
      (X"9F23", X"CF"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"81"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"E7"),
      (X"9F23", X"E7"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"FC"),
      (X"9F23", X"F9"),
      (X"9F23", X"F3"),
      (X"9F23", X"E7"),
      (X"9F23", X"CF"),
      (X"9F23", X"9F"),
      (X"9F23", X"FF"),
      (X"9F23", X"C3"),
      (X"9F23", X"99"),
      (X"9F23", X"91"),
      (X"9F23", X"89"),
      (X"9F23", X"99"),
      (X"9F23", X"99"),
      (X"9F23", X"C3"),
      (X"9F23", X"FF"),
      (X"9F23", X"E7"),
      (X"9F23", X"E7"),
      (X"9F23", X"C7"),
      (X"9F23", X"E7"),
      (X"9F23", X"E7"),
      (X"9F23", X"E7"),
      (X"9F23", X"81"),
      (X"9F23", X"FF"),
      (X"9F23", X"C3"),
      (X"9F23", X"99"),
      (X"9F23", X"F9"),
      (X"9F23", X"F3"),
      (X"9F23", X"CF"),
      (X"9F23", X"9F"),
      (X"9F23", X"81"),
      (X"9F23", X"FF"),
      (X"9F23", X"C3"),
      (X"9F23", X"99"),
      (X"9F23", X"F9"),
      (X"9F23", X"E3"),
      (X"9F23", X"F9"),
      (X"9F23", X"99"),
      (X"9F23", X"C3"),
      (X"9F23", X"FF"),
      (X"9F23", X"F9"),
      (X"9F23", X"F1"),
      (X"9F23", X"E1"),
      (X"9F23", X"99"),
      (X"9F23", X"80"),
      (X"9F23", X"F9"),
      (X"9F23", X"F9"),
      (X"9F23", X"FF"),
      (X"9F23", X"81"),
      (X"9F23", X"9F"),
      (X"9F23", X"83"),
      (X"9F23", X"F9"),
      (X"9F23", X"F9"),
      (X"9F23", X"99"),
      (X"9F23", X"C3"),
      (X"9F23", X"FF"),
      (X"9F23", X"C3"),
      (X"9F23", X"99"),
      (X"9F23", X"9F"),
      (X"9F23", X"83"),
      (X"9F23", X"99"),
      (X"9F23", X"99"),
      (X"9F23", X"C3"),
      (X"9F23", X"FF"),
      (X"9F23", X"81"),
      (X"9F23", X"99"),
      (X"9F23", X"F3"),
      (X"9F23", X"E7"),
      (X"9F23", X"E7"),
      (X"9F23", X"E7"),
      (X"9F23", X"E7"),
      (X"9F23", X"FF"),
      (X"9F23", X"C3"),
      (X"9F23", X"99"),
      (X"9F23", X"99"),
      (X"9F23", X"C3"),
      (X"9F23", X"99"),
      (X"9F23", X"99"),
      (X"9F23", X"C3"),
      (X"9F23", X"FF"),
      (X"9F23", X"C3"),
      (X"9F23", X"99"),
      (X"9F23", X"99"),
      (X"9F23", X"C1"),
      (X"9F23", X"F9"),
      (X"9F23", X"99"),
      (X"9F23", X"C3"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"E7"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"E7"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"E7"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"E7"),
      (X"9F23", X"E7"),
      (X"9F23", X"CF"),
      (X"9F23", X"F1"),
      (X"9F23", X"E7"),
      (X"9F23", X"CF"),
      (X"9F23", X"9F"),
      (X"9F23", X"CF"),
      (X"9F23", X"E7"),
      (X"9F23", X"F1"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"81"),
      (X"9F23", X"FF"),
      (X"9F23", X"81"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"8F"),
      (X"9F23", X"E7"),
      (X"9F23", X"F3"),
      (X"9F23", X"F9"),
      (X"9F23", X"F3"),
      (X"9F23", X"E7"),
      (X"9F23", X"8F"),
      (X"9F23", X"FF"),
      (X"9F23", X"C3"),
      (X"9F23", X"99"),
      (X"9F23", X"F9"),
      (X"9F23", X"F3"),
      (X"9F23", X"E7"),
      (X"9F23", X"FF"),
      (X"9F23", X"E7"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"), -- 0x0FE00
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"F7"),
      (X"9F23", X"E3"),
      (X"9F23", X"C1"),
      (X"9F23", X"80"),
      (X"9F23", X"80"),
      (X"9F23", X"E3"),
      (X"9F23", X"C1"),
      (X"9F23", X"FF"),
      (X"9F23", X"E7"),
      (X"9F23", X"E7"),
      (X"9F23", X"E7"),
      (X"9F23", X"E7"),
      (X"9F23", X"E7"),
      (X"9F23", X"E7"),
      (X"9F23", X"E7"),
      (X"9F23", X"E7"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"CF"),
      (X"9F23", X"CF"),
      (X"9F23", X"CF"),
      (X"9F23", X"CF"),
      (X"9F23", X"CF"),
      (X"9F23", X"CF"),
      (X"9F23", X"CF"),
      (X"9F23", X"CF"),
      (X"9F23", X"F3"),
      (X"9F23", X"F3"),
      (X"9F23", X"F3"),
      (X"9F23", X"F3"),
      (X"9F23", X"F3"),
      (X"9F23", X"F3"),
      (X"9F23", X"F3"),
      (X"9F23", X"F3"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"1F"),
      (X"9F23", X"0F"),
      (X"9F23", X"C7"),
      (X"9F23", X"E7"),
      (X"9F23", X"E7"),
      (X"9F23", X"E7"),
      (X"9F23", X"E7"),
      (X"9F23", X"E3"),
      (X"9F23", X"F0"),
      (X"9F23", X"F8"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"E7"),
      (X"9F23", X"E7"),
      (X"9F23", X"C7"),
      (X"9F23", X"0F"),
      (X"9F23", X"1F"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"3F"),
      (X"9F23", X"3F"),
      (X"9F23", X"3F"),
      (X"9F23", X"3F"),
      (X"9F23", X"3F"),
      (X"9F23", X"3F"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"3F"),
      (X"9F23", X"1F"),
      (X"9F23", X"8F"),
      (X"9F23", X"C7"),
      (X"9F23", X"E3"),
      (X"9F23", X"F1"),
      (X"9F23", X"F8"),
      (X"9F23", X"FC"),
      (X"9F23", X"FC"),
      (X"9F23", X"F8"),
      (X"9F23", X"F1"),
      (X"9F23", X"E3"),
      (X"9F23", X"C7"),
      (X"9F23", X"8F"),
      (X"9F23", X"1F"),
      (X"9F23", X"3F"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"3F"),
      (X"9F23", X"3F"),
      (X"9F23", X"3F"),
      (X"9F23", X"3F"),
      (X"9F23", X"3F"),
      (X"9F23", X"3F"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"FC"),
      (X"9F23", X"FC"),
      (X"9F23", X"FC"),
      (X"9F23", X"FC"),
      (X"9F23", X"FC"),
      (X"9F23", X"FC"),
      (X"9F23", X"FF"),
      (X"9F23", X"C3"),
      (X"9F23", X"81"),
      (X"9F23", X"81"),
      (X"9F23", X"81"),
      (X"9F23", X"81"),
      (X"9F23", X"C3"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"FF"),
      (X"9F23", X"C9"),
      (X"9F23", X"80"),
      (X"9F23", X"80"),
      (X"9F23", X"80"),
      (X"9F23", X"C1"),
      (X"9F23", X"E3"),
      (X"9F23", X"F7"),
      (X"9F23", X"FF"),
      (X"9F23", X"9F"),
      (X"9F23", X"9F"),
      (X"9F23", X"9F"),
      (X"9F23", X"9F"),
      (X"9F23", X"9F"),
      (X"9F23", X"9F"),
      (X"9F23", X"9F"),
      (X"9F23", X"9F"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"F8"),
      (X"9F23", X"F0"),
      (X"9F23", X"E3"),
      (X"9F23", X"E7"),
      (X"9F23", X"E7"),
      (X"9F23", X"3C"),
      (X"9F23", X"18"),
      (X"9F23", X"81"),
      (X"9F23", X"C3"),
      (X"9F23", X"C3"),
      (X"9F23", X"81"),
      (X"9F23", X"18"),
      (X"9F23", X"3C"),
      (X"9F23", X"FF"),
      (X"9F23", X"C3"),
      (X"9F23", X"81"),
      (X"9F23", X"99"),
      (X"9F23", X"99"),
      (X"9F23", X"81"),
      (X"9F23", X"C3"),
      (X"9F23", X"FF"),
      (X"9F23", X"E7"),
      (X"9F23", X"E7"),
      (X"9F23", X"99"),
      (X"9F23", X"99"),
      (X"9F23", X"E7"),
      (X"9F23", X"E7"),
      (X"9F23", X"C3"),
      (X"9F23", X"FF"),
      (X"9F23", X"F9"),
      (X"9F23", X"F9"),
      (X"9F23", X"F9"),
      (X"9F23", X"F9"),
      (X"9F23", X"F9"),
      (X"9F23", X"F9"),
      (X"9F23", X"F9"),
      (X"9F23", X"F9"),
      (X"9F23", X"F7"),
      (X"9F23", X"E3"),
      (X"9F23", X"C1"),
      (X"9F23", X"80"),
      (X"9F23", X"C1"),
      (X"9F23", X"E3"),
      (X"9F23", X"F7"),
      (X"9F23", X"FF"),
      (X"9F23", X"E7"),
      (X"9F23", X"E7"),
      (X"9F23", X"E7"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"E7"),
      (X"9F23", X"E7"),
      (X"9F23", X"E7"),
      (X"9F23", X"3F"),
      (X"9F23", X"3F"),
      (X"9F23", X"CF"),
      (X"9F23", X"CF"),
      (X"9F23", X"3F"),
      (X"9F23", X"3F"),
      (X"9F23", X"CF"),
      (X"9F23", X"CF"),
      (X"9F23", X"E7"),
      (X"9F23", X"E7"),
      (X"9F23", X"E7"),
      (X"9F23", X"E7"),
      (X"9F23", X"E7"),
      (X"9F23", X"E7"),
      (X"9F23", X"E7"),
      (X"9F23", X"E7"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"FC"),
      (X"9F23", X"C1"),
      (X"9F23", X"89"),
      (X"9F23", X"C9"),
      (X"9F23", X"C9"),
      (X"9F23", X"FF"),
      (X"9F23", X"00"),
      (X"9F23", X"80"),
      (X"9F23", X"C0"),
      (X"9F23", X"E0"),
      (X"9F23", X"F0"),
      (X"9F23", X"F8"),
      (X"9F23", X"FC"),
      (X"9F23", X"FE"),
      (X"9F23", X"FF"), -- 0x0FF00
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"0F"),
      (X"9F23", X"0F"),
      (X"9F23", X"0F"),
      (X"9F23", X"0F"),
      (X"9F23", X"0F"),
      (X"9F23", X"0F"),
      (X"9F23", X"0F"),
      (X"9F23", X"0F"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"00"),
      (X"9F23", X"3F"),
      (X"9F23", X"3F"),
      (X"9F23", X"3F"),
      (X"9F23", X"3F"),
      (X"9F23", X"3F"),
      (X"9F23", X"3F"),
      (X"9F23", X"3F"),
      (X"9F23", X"3F"),
      (X"9F23", X"33"),
      (X"9F23", X"33"),
      (X"9F23", X"CC"),
      (X"9F23", X"CC"),
      (X"9F23", X"33"),
      (X"9F23", X"33"),
      (X"9F23", X"CC"),
      (X"9F23", X"CC"),
      (X"9F23", X"FC"),
      (X"9F23", X"FC"),
      (X"9F23", X"FC"),
      (X"9F23", X"FC"),
      (X"9F23", X"FC"),
      (X"9F23", X"FC"),
      (X"9F23", X"FC"),
      (X"9F23", X"FC"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"33"),
      (X"9F23", X"33"),
      (X"9F23", X"CC"),
      (X"9F23", X"CC"),
      (X"9F23", X"00"),
      (X"9F23", X"01"),
      (X"9F23", X"03"),
      (X"9F23", X"07"),
      (X"9F23", X"0F"),
      (X"9F23", X"1F"),
      (X"9F23", X"3F"),
      (X"9F23", X"7F"),
      (X"9F23", X"FC"),
      (X"9F23", X"FC"),
      (X"9F23", X"FC"),
      (X"9F23", X"FC"),
      (X"9F23", X"FC"),
      (X"9F23", X"FC"),
      (X"9F23", X"FC"),
      (X"9F23", X"FC"),
      (X"9F23", X"E7"),
      (X"9F23", X"E7"),
      (X"9F23", X"E7"),
      (X"9F23", X"E0"),
      (X"9F23", X"E0"),
      (X"9F23", X"E7"),
      (X"9F23", X"E7"),
      (X"9F23", X"E7"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"F0"),
      (X"9F23", X"F0"),
      (X"9F23", X"F0"),
      (X"9F23", X"F0"),
      (X"9F23", X"E7"),
      (X"9F23", X"E7"),
      (X"9F23", X"E7"),
      (X"9F23", X"E0"),
      (X"9F23", X"E0"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"07"),
      (X"9F23", X"07"),
      (X"9F23", X"E7"),
      (X"9F23", X"E7"),
      (X"9F23", X"E7"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"E0"),
      (X"9F23", X"E0"),
      (X"9F23", X"E7"),
      (X"9F23", X"E7"),
      (X"9F23", X"E7"),
      (X"9F23", X"E7"),
      (X"9F23", X"E7"),
      (X"9F23", X"E7"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"E7"),
      (X"9F23", X"E7"),
      (X"9F23", X"E7"),
      (X"9F23", X"E7"),
      (X"9F23", X"E7"),
      (X"9F23", X"E7"),
      (X"9F23", X"07"),
      (X"9F23", X"07"),
      (X"9F23", X"E7"),
      (X"9F23", X"E7"),
      (X"9F23", X"E7"),
      (X"9F23", X"3F"),
      (X"9F23", X"3F"),
      (X"9F23", X"3F"),
      (X"9F23", X"3F"),
      (X"9F23", X"3F"),
      (X"9F23", X"3F"),
      (X"9F23", X"3F"),
      (X"9F23", X"3F"),
      (X"9F23", X"1F"),
      (X"9F23", X"1F"),
      (X"9F23", X"1F"),
      (X"9F23", X"1F"),
      (X"9F23", X"1F"),
      (X"9F23", X"1F"),
      (X"9F23", X"1F"),
      (X"9F23", X"1F"),
      (X"9F23", X"F8"),
      (X"9F23", X"F8"),
      (X"9F23", X"F8"),
      (X"9F23", X"F8"),
      (X"9F23", X"F8"),
      (X"9F23", X"F8"),
      (X"9F23", X"F8"),
      (X"9F23", X"F8"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"FC"),
      (X"9F23", X"FC"),
      (X"9F23", X"FC"),
      (X"9F23", X"FC"),
      (X"9F23", X"FC"),
      (X"9F23", X"FC"),
      (X"9F23", X"00"),
      (X"9F23", X"00"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"0F"),
      (X"9F23", X"0F"),
      (X"9F23", X"0F"),
      (X"9F23", X"0F"),
      (X"9F23", X"F0"),
      (X"9F23", X"F0"),
      (X"9F23", X"F0"),
      (X"9F23", X"F0"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"E7"),
      (X"9F23", X"E7"),
      (X"9F23", X"E7"),
      (X"9F23", X"07"),
      (X"9F23", X"07"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"0F"),
      (X"9F23", X"0F"),
      (X"9F23", X"0F"),
      (X"9F23", X"0F"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"FF"),
      (X"9F23", X"0F"),
      (X"9F23", X"0F"),
      (X"9F23", X"0F"),
      (X"9F23", X"0F"),
      (X"9F23", X"F0"),
      (X"9F23", X"F0"),
      (X"9F23", X"F0"),
      (X"9F23", X"F0")
   );

   signal wr_index : integer := 0;

begin

   -- This is a temporary process that populates the VRAM
   p_wr : process (clk_i)
   begin
      if rising_edge(clk_i) then
         wr_en_o <= '0';
         if wr_index < wr_default'length then
            wr_addr_o <= wr_default(wr_index).addr(2 downto 0);
            wr_en_o   <= '1';
            wr_data_o <= wr_default(wr_index).data;
            wr_index  <= wr_index + 1;
         end if;
      end if;
   end process p_wr;

end architecture structural;


--------------------------------------
-- The Control Logic
--
-- This uses a ROM containing up to eight microcodes for each instruction.

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.std_logic_arith.all;

entity ctl is
   port (
      clk_i  : in  std_logic;
      rst_i  : in  std_logic;
      irq_i  : in  std_logic;
      data_i : in  std_logic_vector( 7 downto 0);

      mem_rden_o      : out std_logic;                      -- Read from memory
      mem_wren_o      : out std_logic;                      -- Write to memory
      mem_addr_wren_o : out std_logic_vector(1 downto 0);   -- Write to address hold register
      mem_addr_sel_o  : out std_logic_vector(3 downto 0);   -- Memory address select
      mem_data_sel_o  : out std_logic_vector(1 downto 0);   -- Memory data select
      reg_wren_o      : out std_logic;                      -- Write to register file
      reg_nr_o        : out std_logic_vector(1 downto 0);   -- Register number
      pc_sel_o        : out std_logic_vector(1 downto 0);   -- PC relect
      sp_sel_o        : out std_logic_vector(1 downto 0);   -- Stack pointer update
      alu_func_o      : out std_logic_vector(3 downto 0);   -- ALU function
      clc_o           : out std_logic;                      -- Clear carry
      sr_alu_wren_o   : out std_logic;                      -- Write status register
      irq_mask_wr_o   : out std_logic_vector(1 downto 0);   -- Write to irq mask bit

      debug_o : out std_logic_vector(10 downto 0)
   );
end ctl;

architecture Structural of ctl is

   signal cnt_r   : std_logic_vector(2 downto 0) := (others => '0');
   signal inst_r  : std_logic_vector(7 downto 0) := (others => '0');
   signal last    : std_logic;
   signal invalid : std_logic;

   signal ctl     : std_logic_vector(26 downto 0);
   signal irq_l   : std_logic := '0';
   signal rst_l   : std_logic := '0';

   subtype micro_op_type is std_logic_vector(26 downto 0);
   type micro_op_rom_type is array(0 to 8*256-1) of micro_op_type;

   constant C_READ_NEXT_BYTE : micro_op_type :=
      B"00_0_0_0_0_0000_00_00_00_0_00_0000_00_0_1";

   constant C_NOT_IMPLEMENTED : micro_op_type := 
      B"00_1_0_0_0_0000_00_00_00_0_00_0000_00_0_0";

   constant micro_op_rom : micro_op_rom_type := (
   -- 00 BRK b
            C_READ_NEXT_BYTE,
            B"00_0_0_0_0_0000_10_11_00_0_01_0010_00_1_0",
            B"00_0_0_0_0_0000_10_11_00_0_10_0010_00_1_0",
            B"11_0_0_0_0_0000_10_11_00_0_11_0010_00_1_0",
            B"00_0_0_0_0_0000_00_11_00_0_00_1000_01_0_1",
            B"00_0_1_0_0_0000_00_01_00_0_00_1001_10_0_1",
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- 01 ORA (d,X)
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- 02
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- 03
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- 04
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- 05 ORA d
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- 06 ASL d
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- 07
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- 08 PHP
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- 09 ORA #
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- 0A ASL A
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- 0B
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- 0C
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- 0D ORA a
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- 0E ASL a
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- 0F
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   --
   -- 10 BPL r
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- 11 ORA (d),Y
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- 12
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- 13
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- 14
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- 15 ORA d,X
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- 16 ASL d,X
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- 17
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- 18 CLC
            C_READ_NEXT_BYTE,
            B"00_0_1_0_1_0000_00_11_00_0_00_0000_00_0_0",
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- 19 ORA a,Y
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- 1A
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- 1B
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- 1C
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- 1D ORA a,X
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- 1E ASL a,X
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- 1F
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   --
   -- 20 JSR a
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- 21 AND (d,X)
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- 22
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- 23
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- 24 BIT d
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- 25 AND d
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- 26 ROL d
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- 27
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- 28 PLP
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- 29 AND #
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- 2A ROL A
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- 2B
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- 2C BIT a
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- 2D AND a
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- 2E ROL a
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- 2F
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   --
   -- 30 BMI r
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- 31 AND (d),Y
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- 32
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- 33
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- 34
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- 35 AND d,X
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- 36 ROL d,X
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- 37
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- 38 SEC
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- 39 AND a,Y
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- 3A
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- 3B
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- 3C
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- 3D AND a,X
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- 3E ROL a,X
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- 3F
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   --
   -- 40 RTI
            C_READ_NEXT_BYTE,
            B"00_0_0_0_0_0000_01_11_00_0_00_0000_00_0_0",
            B"01_0_0_0_0_0000_01_11_00_0_00_0010_00_0_1",
            B"00_0_0_0_0_0000_01_11_00_0_00_0010_01_0_1",
            B"00_0_1_0_0_0000_00_01_00_0_00_0010_00_0_1",
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- 41 EOR (d,X)
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- 42
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- 43
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- 44
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- 45 EOR d
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- 46 LSR d
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- 47
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- 48 PHA
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- 49 EOR #
            C_READ_NEXT_BYTE,
            B"00_0_1_1_0_0010_00_00_00_1_00_0000_00_0_1",
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- 4A LSR A
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- 4B
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- 4C JMP a
            C_READ_NEXT_BYTE,
            B"00_0_0_0_0_0000_00_00_00_0_00_0000_01_0_1",
            B"00_0_1_0_0_0000_00_01_00_0_00_0000_00_0_1",
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- 4D EOR a
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- 4E LSR a
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- 4F
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   --
   -- 50 BVC r
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- 51 EOR (d),Y
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- 52
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- 53
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- 54
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- 55 EOR d,X
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- 56 LSR d,X
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- 57
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- 58 CLI
            C_READ_NEXT_BYTE,
            B"10_0_1_0_0_0000_00_11_00_0_00_0000_00_0_0",
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- 59 EOR a,Y
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- 5A
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- 5B
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- 5C
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- 5D EOR a,X
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- 5E LSR a,X
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- 5F
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   --
   -- 60 RTS
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- 61 ADC (d,X)
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- 62
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- 63
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- 64
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- 65 ADC d
            C_READ_NEXT_BYTE,
            B"00_0_0_0_0_0000_00_00_00_0_00_0000_01_0_1",
            B"00_0_1_1_0_0011_00_11_00_1_00_0001_00_0_1",
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- 66 ROR d
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- 67
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- 68 PLA
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- 69 ADC #
            C_READ_NEXT_BYTE,
            B"00_0_1_1_0_0011_00_00_00_1_00_0000_00_0_1",
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- 6A ROR A
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- 6B
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- 6C JMP (a)
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- 6D ADC a
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- 6E ROR a
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- 6F
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   --
   -- 70 BVS r
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- 71 ADC (d),Y
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- 72
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- 73
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- 74
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- 75 ADC d,X
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- 76 ROR d,X
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- 77
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- 78 SEI
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- 79 ADC a,Y
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- 7A
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- 7B
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- 7C
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- 7D ADC a,X
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- 7E ROR a,X
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- 7F
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   --
   -- 80
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- 81 STA (d,X)
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- 82
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- 83
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- 84 STY
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- 85 STA d
            C_READ_NEXT_BYTE,
            B"00_0_0_0_0_0000_00_00_00_0_00_0000_01_0_1",
            B"00_0_1_0_0_0000_00_11_00_0_00_0001_00_1_0",
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- 86 STX d
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- 87
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- 88 DEY
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- 89
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- 8A TXA
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- 8B
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- 8C STY a
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- 8D STA a
            C_READ_NEXT_BYTE,
            B"00_0_0_0_0_0000_00_00_00_0_00_0000_01_0_1",
            B"00_0_0_0_0_0000_00_00_00_0_00_0000_10_0_1",
            B"00_0_1_0_0_0000_00_11_00_0_00_0011_00_1_0",
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- 8E STX a
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- 8F
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   --
   -- 90 BCC r
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- 91 STA (d),Y
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- 92
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- 93
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- 94 STY d,X
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- 95 STA d,X
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- 96 STX d,Y
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- 97
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- 98 TYA
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- 99 STA a,Y
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- 9A TXS
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- 9B
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- 9C
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- 9D STA a,X
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- 9E
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- 9F
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   --
   -- A0 LDY #
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- A1 LDA (d,X)
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- A2 LDX #
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- A3
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- A4 LDY d
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- A5 LDA d
            C_READ_NEXT_BYTE,
            B"00_0_0_0_0_0000_00_00_00_0_00_0000_01_0_1",
            B"00_0_1_0_0_0101_00_11_00_1_00_0001_00_0_1",
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- A6 LDX d
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- A7
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- A8 TAY
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- A9 LDA #
            C_READ_NEXT_BYTE,
            B"00_0_1_0_0_0101_00_00_00_1_00_0000_00_0_1",
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- AA TAX
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- AB
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- AC LDY a
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- AD LDA a
            C_READ_NEXT_BYTE,
            B"00_0_0_0_0_0000_00_00_00_0_00_0000_01_0_1",
            B"00_0_0_0_0_0000_00_00_00_0_00_0000_10_0_1",
            B"00_0_1_0_0_0101_00_11_00_1_00_0011_00_0_1",
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- AE LDX a
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- AF
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   --
   -- B0 BCS r
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- B1 LDA (d),Y
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- B2
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- B3
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- B4 LDY d,X
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- B5 LDA d,X
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- B6 LDX d,Y
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- B7
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- B8 CLV
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- B9 LDA a,Y
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- BA TSX
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- BB
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- BC LDY a,X
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- BD LDA a,X
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- BE LDX a,Y
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- BF
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   --
   -- C0 CPY #
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- C1 CMP (d,X)
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- C2
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- C3
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- C4 CPY d
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- C5 CMP d
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- C6 DEC d
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- C7
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- C8 INY
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- C9 CMP #
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- CA DEX
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- CB
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- CC CPY a
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- CD CMP a
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- CE DEC a
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- CF
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   --
   -- D0 BNE r
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- D1 CMP (d),Y
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- D2
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- D3
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- D4
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- D5 CMP d,X
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- D6 DEC d,X
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- D7
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- D8 CLD
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- D9 CMP a,Y
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- DA
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- DB
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- DC
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- DD CMP a,X
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- DE DEC a,X
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- DF
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   --
   -- E0 CPX #
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- E1 SBC (d,X)
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- E2
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- E3
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- E4 CPX d
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- E5 SBC d
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- E6 INC d
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- E7
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- E8 INX
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- E9 SBC #
            C_READ_NEXT_BYTE,
            B"00_0_1_1_0_0111_00_00_00_1_00_0000_00_0_1",
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- EA NOP
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- EB
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- EC CPX a
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- ED SBC a
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- EE INC a
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- EF
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   --
   -- F0 BEQ r
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- F1 SBC (d),Y
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- F2
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- F3
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- F4
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- F5 SBC d,X
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- F6 INC d,X
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- F7
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- F8 SED
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- F9 SBC a,Y
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- FA
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- FB
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- FC
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- FD SBC a,X
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- FE INC a,X
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
   -- FF
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED,
            C_NOT_IMPLEMENTED
         );

begin

   -- Check for illegal or unimplemented instructions.
   p_assert : process (clk_i)
   begin 
      if rising_edge(clk_i) then
         if rst_i = '0' then
            assert invalid = '0' report "Invalid opcode" severity failure;
         end if;
      end if;
   end process p_assert;


   -- Store the microinstruction counter
   p_cnt : process (clk_i)
   begin
      if rising_edge(clk_i) then
         cnt_r <= cnt_r + 1;

         if last = '1' then
            cnt_r <= (others => '0');

            if irq_i = '1' then
               cnt_r <= "001";
            end if;
         end if;

         if rst_i = '1' then
            cnt_r <= "011";
         end if;
      end if;
   end process p_cnt;


   -- Store the current instruction
   p_inst : process (clk_i)
   begin
      if rising_edge(clk_i) then
         if cnt_r = 0 then
            inst_r <= data_i;
         end if;

         if last = '1' and irq_i = '1' then
            inst_r <= X"00";
         end if;

         if rst_i = '1' then
            inst_r <= X"00";
         end if;
      end if;
   end process p_inst;


   -- Latch reset and interrupt
   p_irq_reset : process (clk_i)
   begin
      if rising_edge(clk_i) then
         if last = '1' then
            irq_l <= irq_i;
            rst_l <= irq_i;
         end if;

         if rst_i = '1' then
            irq_l <= '0';
            rst_l <= rst_i;
         end if;
      end if;
   end process p_irq_reset;

   -- Combinatorial process
   process (cnt_r, inst_r)
   begin
      ctl <= micro_op_rom(conv_integer(inst_r & cnt_r));
   end process;

   -- Drive output signals
   mem_rden_o      <= ctl(0);
   mem_wren_o      <= ctl(1);
   mem_addr_wren_o <= ctl(3 downto 2);
   mem_addr_sel_o  <= ctl(7 downto 4) when ctl(7) = '0'
                      else '1' & rst_l & irq_l & ctl(4);
   mem_data_sel_o  <= ctl(9 downto 8);
   reg_wren_o      <= ctl(10);
   reg_nr_o        <= ctl(12 downto 11);
   pc_sel_o        <= ctl(14 downto 13);
   sp_sel_o        <= ctl(16 downto 15);
   alu_func_o      <= ctl(20 downto 17);
   clc_o           <= ctl(21);
   sr_alu_wren_o   <= ctl(22);
   last            <= ctl(23);
   invalid         <= ctl(24);
   irq_mask_wr_o   <= ctl(26 downto 25);

   debug_o( 7 downto 0) <= inst_r;
   debug_o(10 downto 8) <= cnt_r;

end architecture Structural;



   -- Default palette. Mapping from 8-bits to 12-bits.
   -- Copied from x16-emulator.
   X"000", X"fff", X"800", X"afe", X"c4c", X"0c5", X"00a", X"ee7", X"d85", X"640", X"f77", X"333", X"777", X"af6", X"08f", X"bbb",
   X"000", X"111", X"222", X"333", X"444", X"555", X"666", X"777", X"888", X"999", X"aaa", X"bbb", X"ccc", X"ddd", X"eee", X"fff",
   X"211", X"433", X"644", X"866", X"a88", X"c99", X"fbb", X"211", X"422", X"633", X"844", X"a55", X"c66", X"f77", X"200", X"411",
   X"611", X"822", X"a22", X"c33", X"f33", X"200", X"400", X"600", X"800", X"a00", X"c00", X"f00", X"221", X"443", X"664", X"886",
   X"aa8", X"cc9", X"feb", X"211", X"432", X"653", X"874", X"a95", X"cb6", X"fd7", X"210", X"431", X"651", X"862", X"a82", X"ca3",
   X"fc3", X"210", X"430", X"640", X"860", X"a80", X"c90", X"fb0", X"121", X"343", X"564", X"786", X"9a8", X"bc9", X"dfb", X"121",
   X"342", X"463", X"684", X"8a5", X"9c6", X"bf7", X"120", X"241", X"461", X"582", X"6a2", X"8c3", X"9f3", X"120", X"240", X"360",
   X"480", X"5a0", X"6c0", X"7f0", X"121", X"343", X"465", X"686", X"8a8", X"9ca", X"bfc", X"121", X"242", X"364", X"485", X"5a6",
   X"6c8", X"7f9", X"020", X"141", X"162", X"283", X"2a4", X"3c5", X"3f6", X"020", X"041", X"061", X"082", X"0a2", X"0c3", X"0f3",
   X"122", X"344", X"466", X"688", X"8aa", X"9cc", X"bff", X"122", X"244", X"366", X"488", X"5aa", X"6cc", X"7ff", X"022", X"144",
   X"166", X"288", X"2aa", X"3cc", X"3ff", X"022", X"044", X"066", X"088", X"0aa", X"0cc", X"0ff", X"112", X"334", X"456", X"668",
   X"88a", X"9ac", X"bcf", X"112", X"224", X"346", X"458", X"56a", X"68c", X"79f", X"002", X"114", X"126", X"238", X"24a", X"35c",
   X"36f", X"002", X"014", X"016", X"028", X"02a", X"03c", X"03f", X"112", X"334", X"546", X"768", X"98a", X"b9c", X"dbf", X"112",
   X"324", X"436", X"648", X"85a", X"96c", X"b7f", X"102", X"214", X"416", X"528", X"62a", X"83c", X"93f", X"102", X"204", X"306",
   X"408", X"50a", X"60c", X"70f", X"212", X"434", X"646", X"868", X"a8a", X"c9c", X"fbe", X"211", X"423", X"635", X"847", X"a59",
   X"c6b", X"f7d", X"201", X"413", X"615", X"826", X"a28", X"c3a", X"f3c", X"201", X"403", X"604", X"806", X"a08", X"c09", X"f0b",


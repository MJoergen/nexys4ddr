library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

package vga_bitmap_pkg is

   -- These are the pixel dimensions of each character.
   -- It is a monospace font, for simplicity. Non-monospace is too hard :-)
   constant CHAR_WIDTH  : integer := 11;
   constant CHAR_HEIGHT : integer := 16;

   subtype vga_bitmap_t is std_logic_vector(0 to CHAR_WIDTH * CHAR_HEIGHT - 1);

   constant vga_bitmap_char_0 : vga_bitmap_t := (
      "00000000000" &
      "00000000000" &
      "00001110000" &
      "00010001000" &
      "00100000100" &
      "00100000100" &
      "00100000100" &
      "00100000100" &
      "00100000100" &
      "00100000100" &
      "00100000100" &
      "00100000100" &
      "00010001000" &
      "00001110000" &
      "00000000000" &
      "00000000000");

   constant vga_bitmap_char_1 : vga_bitmap_t := (
      "00000000000" &
      "00000000000" &
      "00001100000" &
      "00110100000" &
      "00000100000" &
      "00000100000" &
      "00000100000" &
      "00000100000" &
      "00000100000" &
      "00000100000" &
      "00000100000" &
      "00000100000" &
      "00000100000" &
      "00111111100" &
      "00000000000" &
      "00000000000");

   constant vga_bitmap_char_2 : vga_bitmap_t := (
      "00000000000" &
      "00000000000" &
      "00001110000" &
      "00010001000" &
      "00100000100" &
      "00000000100" &
      "00000000100" &
      "00000001000" &
      "00000010000" &
      "00000100000" &
      "00001000000" &
      "00010000000" &
      "00100000000" &
      "00111111100" &
      "00000000000" &
      "00000000000");

   constant vga_bitmap_char_3 : vga_bitmap_t := (
      "00000000000" &
      "00000000000" &
      "00001110000" &
      "00010001000" &
      "00100000100" &
      "00000000100" &
      "00000001000" &
      "00000110000" &
      "00000001000" &
      "00000000100" &
      "00000000100" &
      "00100000100" &
      "00010001000" &
      "00001110000" &
      "00000000000" &
      "00000000000");

   constant vga_bitmap_char_4 : vga_bitmap_t := (
      "00000000000" &
      "00000000000" &
      "00000001000" &
      "00000011000" &
      "00000101000" &
      "00001001000" &
      "00010001000" &
      "00111111100" &
      "00000001000" &
      "00000001000" &
      "00000001000" &
      "00000001000" &
      "00000001000" &
      "00000001000" &
      "00000000000" &
      "00000000000");

   constant vga_bitmap_char_5 : vga_bitmap_t := (
      "00000000000" &
      "00000000000" &
      "00111111100" &
      "00100000000" &
      "00100000000" &
      "00100000000" &
      "00100000000" &
      "00111110000" &
      "00000001000" &
      "00000000100" &
      "00000000100" &
      "00100000100" &
      "00010001000" &
      "00001110000" &
      "00000000000" &
      "00000000000");

   constant vga_bitmap_char_6 : vga_bitmap_t := (
      "00000000000" &
      "00000000000" &
      "00001111000" &
      "00010000000" &
      "00100000000" &
      "00100000000" &
      "00100000000" &
      "00111110000" &
      "00110001000" &
      "00100000100" &
      "00100000100" &
      "00100000100" &
      "00010001000" &
      "00001110000" &
      "00000000000" &
      "00000000000");

   constant vga_bitmap_char_7 : vga_bitmap_t := (
      "00000000000" &
      "00000000000" &
      "00111111100" &
      "00000000100" &
      "00000000100" &
      "00000001000" &
      "00000001000" &
      "00000010000" &
      "00000010000" &
      "00000100000" &
      "00000100000" &
      "00001000000" &
      "00001000000" &
      "00001000000" &
      "00000000000" &
      "00000000000");

   constant vga_bitmap_char_8 : vga_bitmap_t := (
      "00000000000" &
      "00000000000" &
      "00001110000" &
      "00010001000" &
      "00100000100" &
      "00100000100" &
      "00010001000" &
      "00001110000" &
      "00010001000" &
      "00100000100" &
      "00100000100" &
      "00100000100" &
      "00010001000" &
      "00001110000" &
      "00000000000" &
      "00000000000");

   constant vga_bitmap_char_9 : vga_bitmap_t := (
      "00000000000" &
      "00000000000" &
      "00001110000" &
      "00010001000" &
      "00100000100" &
      "00100000100" &
      "00100000100" &
      "00010000100" &
      "00001111100" &
      "00000000100" &
      "00000000100" &
      "00000000100" &
      "00100001000" &
      "00011110000" &
      "00000000000" &
      "00000000000");

   constant vga_bitmap_char_A : vga_bitmap_t := (
      "00000000000" &
      "00000000000" &
      "00001110000" &
      "00010001000" &
      "00010001000" &
      "00010001000" &
      "00010001000" &
      "00010001000" &
      "00111111100" &
      "00100000100" &
      "00100000100" &
      "00100000100" &
      "00100000100" &
      "00100000100" &
      "00000000000" &
      "00000000000");

   constant vga_bitmap_char_B : vga_bitmap_t := (
      "00000000000" &
      "00000000000" &
      "00111110000" &
      "00100001000" &
      "00100000100" &
      "00100000100" &
      "00100001000" &
      "00111110000" &
      "00100001000" &
      "00100000100" &
      "00100000100" &
      "00100000100" &
      "00100001000" &
      "00111110000" &
      "00000000000" &
      "00000000000");

   constant vga_bitmap_char_C : vga_bitmap_t := (
      "00000000000" &
      "00000000000" &
      "00001111000" &
      "00010000100" &
      "00100000000" &
      "00100000000" &
      "00100000000" &
      "00100000000" &
      "00100000000" &
      "00100000000" &
      "00100000000" &
      "00100000000" &
      "00010000100" &
      "00001111000" &
      "00000000000" &
      "00000000000");

   constant vga_bitmap_char_D : vga_bitmap_t := (
      "00000000000" &
      "00000000000" &
      "00111110000" &
      "00100001000" &
      "00100000100" &
      "00100000100" &
      "00100000100" &
      "00100000100" &
      "00100000100" &
      "00100000100" &
      "00100000100" &
      "00100000100" &
      "00100001000" &
      "00111110000" &
      "00000000000" &
      "00000000000");

   constant vga_bitmap_char_E : vga_bitmap_t := (
      "00000000000" &
      "00000000000" &
      "00111111100" &
      "00100000000" &
      "00100000000" &
      "00100000000" &
      "00100000000" &
      "00111111000" &
      "00100000000" &
      "00100000000" &
      "00100000000" &
      "00100000000" &
      "00100000000" &
      "00111111100" &
      "00000000000" &
      "00000000000");

   constant vga_bitmap_char_F : vga_bitmap_t := (
      "00000000000" &
      "00000000000" &
      "00111111100" &
      "00100000000" &
      "00100000000" &
      "00100000000" &
      "00100000000" &
      "00111111000" &
      "00100000000" &
      "00100000000" &
      "00100000000" &
      "00100000000" &
      "00100000000" &
      "00100000000" &
      "00000000000" &
      "00000000000");

   -- TBD: Do the rest of the alphabet.

   type vga_letters_t is array (0 to 15) of vga_bitmap_t;

   constant vga_letters : vga_letters_t := (
      vga_bitmap_char_0,
      vga_bitmap_char_1,
      vga_bitmap_char_2,
      vga_bitmap_char_3,
      vga_bitmap_char_4,
      vga_bitmap_char_5,
      vga_bitmap_char_6,
      vga_bitmap_char_7,
      vga_bitmap_char_8,
      vga_bitmap_char_9,
      vga_bitmap_char_A,
      vga_bitmap_char_B,
      vga_bitmap_char_C,
      vga_bitmap_char_D,
      vga_bitmap_char_E,
      vga_bitmap_char_F);

   -- Define some common colours
   constant vga_white   : std_logic_vector(11 downto 0) := "1111" & "1111" & "1111";
   constant vga_light   : std_logic_vector(11 downto 0) := "1100" & "1100" & "1100";
   constant vga_gray    : std_logic_vector(11 downto 0) := "1000" & "1000" & "1000";
   constant vga_dark    : std_logic_vector(11 downto 0) := "0100" & "0100" & "0100";
   constant vga_black   : std_logic_vector(11 downto 0) := "0000" & "0000" & "0000";
   constant vga_red     : std_logic_vector(11 downto 0) := "1111" & "0000" & "0000";
   constant vga_green   : std_logic_vector(11 downto 0) := "0000" & "1111" & "0000";
   constant vga_blue    : std_logic_vector(11 downto 0) := "0000" & "0000" & "1111";
   constant vga_cyan    : std_logic_vector(11 downto 0) := "0000" & "1111" & "1111";
   constant vga_magenta : std_logic_vector(11 downto 0) := "1111" & "0000" & "1111";
   constant vga_yellow  : std_logic_vector(11 downto 0) := "1111" & "1111" & "0000";

end package vga_bitmap_pkg;


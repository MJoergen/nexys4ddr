library ieee;
use ieee.std_logic_1164.all;

-- This block is a dummy block that generates a number of writes from the CPU,
-- simulating the KERNAL/BASIC ROM.
-- It is also used during simulation to test the VERA block.
--
-- Upon startup the KERNAL/BASIC performs the following sequence of writes to the VERA:
-- 1. 0x0F800 - 0x0FFFF : Tile data.
-- 2. 0xF3000 - 0xF3009 : Layer 2.  Values 01:06:00:00:00:3E:00:00:00:00
-- 3. 0xF0000 - 0xF0008 : Composer. Values 01:80:80:0E:00:80:00:E0:28
-- 4. 0x00000 - 0x03FFF : Clear screen. Values 20:61 repeated.
-- 5. 0x00000 - 0x008FF : Display welcome screen.
--
-- The default values of the composer settings are interpreted as follows:
-- * VGA output
-- * HSCALE = VSCALE = 0x80, which means 1 output pixel for every input pixel.
-- * HSTART = 0, HSTOP = 640
-- * VSTART = 0, VSTOP = 480
-- 
-- The default values of the layer settings are interpreted as follows:
-- * MODE = 0, which means 16 colour text mode
-- * MAPW = 2, which means 128 tiles wide
-- * MAPH = 1, which means 64 tiles high
-- * TILEW = TILEH = 0, which means each tile is 8x8
-- * MAPBASE = 0, which means the MAP area starts at 0x00000
-- * TILEBASE = 0x3E00, which means the TILE area starts at 0x0F800
-- * HSCROLL = VSCROLL = 0

entity cpu_dummy is
   port (
      clk_i     : in  std_logic;
      addr_o    : out std_logic_vector(2 downto 0);
      wr_en_o   : out std_logic;
      wr_data_o : out std_logic_vector(7 downto 0);
      rd_en_o   : out std_logic;
      rd_data_i : in  std_logic_vector(7 downto 0)
   );
end cpu_dummy;

architecture structural of cpu_dummy is

   signal exp_data_r : std_logic_vector(7 downto 0);

   -- This defines a type containing an array of bytes
   type command is record
      addr  : std_logic_vector(15 downto 0);
      data  : std_logic_vector( 7 downto 0);
      wr_en : std_logic;
   end record command;
   type command_vector is array (natural range <>) of command;

   constant commands : command_vector := (
      -- Configure layer 1
      (X"9F25", X"00", '1'), -- Select address port 0
      (X"9F20", X"00", '1'),
      (X"9F21", X"30", '1'),
      (X"9F22", X"1F", '1'), -- Set address to 0xF3000 and increment to 1.
      (X"9F23", X"01", '1'), -- 0xF3000
      (X"9F23", X"06", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"3E", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),

      (X"9F20", X"0A", '0'), -- VERIFY read from address 0x9F20
      (X"9F21", X"30", '0'), -- VERIFY read from address 0x9F21
      (X"9F22", X"1F", '0'), -- VERIFY read from address 0x9F22

      (X"9F20", X"04", '1'),
      (X"9F21", X"30", '1'),
      (X"9F22", X"1F", '1'), -- Set address to 0xF3004 and increment to 1.
      (X"9F23", X"00", '0'), -- VERIFY read from configuraton register 0xF3004
      (X"9F23", X"3E", '0'), -- VERIFY read from configuraton register 0xF3005

      (X"9F20", X"06", '1'),
      (X"9F21", X"10", '1'),
      (X"9F22", X"1F", '1'), -- Set address to 0xF1003 and increment to 1.
      (X"9F23", X"FE", '0'), -- VERIFY read from configuraton register 0xF1006
      (X"9F23", X"0A", '0'), -- VERIFY read from configuraton register 0xF1007

      -- Configure display composer
      (X"9F20", X"00", '1'),
      (X"9F21", X"00", '1'),
      (X"9F22", X"1F", '1'), -- Set address to 0xF0000 and increment to 1.
      (X"9F23", X"01", '1'), -- 0xF0000
      (X"9F23", X"80", '1'),
      (X"9F23", X"80", '1'),
      (X"9F23", X"0E", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"80", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"E0", '1'),
      (X"9F23", X"28", '1'),

      -- The first part is the map area, i.e. the characters and colours.
      (X"9F20", X"00", '1'),
      (X"9F21", X"00", '1'),
      (X"9F22", X"10", '1'), -- Set address to 0x00000 and increment to 1.
      (X"9F23", X"5F", '1'), -- 0x00000
      (X"9F23", X"64", '1'),
      (X"9F23", X"A0", '1'),
      (X"9F23", X"64", '1'),
      (X"9F23", X"A0", '1'),
      (X"9F23", X"64", '1'),
      (X"9F23", X"DF", '1'),
      (X"9F23", X"64", '1'),
      (X"9F23", X"20", '1'),
      (X"9F23", X"64", '1'),
      (X"9F23", X"20", '1'),
      (X"9F23", X"64", '1'),
      (X"9F23", X"20", '1'),
      (X"9F23", X"64", '1'),
      (X"9F23", X"E9", '1'),
      (X"9F23", X"64", '1'),
      (X"9F23", X"A0", '1'), -- 0x00010
      (X"9F23", X"64", '1'),
      (X"9F23", X"A0", '1'),
      (X"9F23", X"64", '1'),
      (X"9F23", X"69", '1'),
      (X"9F23", X"64", '1'),

      (X"9F20", X"02", '1'),
      (X"9F21", X"00", '1'),
      (X"9F22", X"10", '1'), -- Set address to 0x00002 and increment to 1.
      (X"9F23", X"A0", '0'), -- VERIFY read from VRAM address 0x00002
      (X"9F23", X"64", '0'), -- VERIFY read from VRAM address 0x00003

      (X"9F20", X"00", '1'),
      (X"9F21", X"01", '1'), -- Set address to 0x00100
      (X"9F23", X"20", '1'), -- 0x00100
      (X"9F23", X"6E", '1'),
      (X"9F23", X"5F", '1'),
      (X"9F23", X"6E", '1'),
      (X"9F23", X"A0", '1'),
      (X"9F23", X"6E", '1'),
      (X"9F23", X"A0", '1'),
      (X"9F23", X"6E", '1'),
      (X"9F23", X"DF", '1'),
      (X"9F23", X"6E", '1'),
      (X"9F23", X"20", '1'),
      (X"9F23", X"6E", '1'),
      (X"9F23", X"E9", '1'),
      (X"9F23", X"6E", '1'),
      (X"9F23", X"A0", '1'),
      (X"9F23", X"6E", '1'),
      (X"9F23", X"A0", '1'), -- 0x00110
      (X"9F23", X"6E", '1'),
      (X"9F23", X"69", '1'),
      (X"9F23", X"6E", '1'),
      (X"9F23", X"20", '1'),
      (X"9F23", X"61", '1'),
      (X"9F23", X"20", '1'),
      (X"9F23", X"61", '1'),
      (X"9F23", X"2A", '1'),
      (X"9F23", X"61", '1'),
      (X"9F23", X"2A", '1'),
      (X"9F23", X"61", '1'),
      (X"9F23", X"2A", '1'),
      (X"9F23", X"61", '1'),
      (X"9F23", X"2A", '1'),
      (X"9F23", X"61", '1'),
      (X"9F23", X"20", '1'), -- 0x00120
      (X"9F23", X"61", '1'),
      (X"9F23", X"03", '1'),
      (X"9F23", X"61", '1'),
      (X"9F23", X"0F", '1'),
      (X"9F23", X"61", '1'),
      (X"9F23", X"0D", '1'),
      (X"9F23", X"61", '1'),
      (X"9F23", X"0D", '1'),
      (X"9F23", X"61", '1'),
      (X"9F23", X"01", '1'),
      (X"9F23", X"61", '1'),
      (X"9F23", X"0E", '1'),
      (X"9F23", X"61", '1'),
      (X"9F23", X"04", '1'),
      (X"9F23", X"61", '1'),
      (X"9F23", X"05", '1'), -- 0x00130
      (X"9F23", X"61", '1'),
      (X"9F23", X"12", '1'),
      (X"9F23", X"61", '1'),
      (X"9F23", X"20", '1'),
      (X"9F23", X"61", '1'),
      (X"9F23", X"18", '1'),
      (X"9F23", X"61", '1'),
      (X"9F23", X"31", '1'),
      (X"9F23", X"61", '1'),
      (X"9F23", X"36", '1'),
      (X"9F23", X"61", '1'),
      (X"9F23", X"20", '1'),
      (X"9F23", X"61", '1'),
      (X"9F23", X"02", '1'),
      (X"9F23", X"61", '1'),
      (X"9F23", X"01", '1'), -- 0x00140
      (X"9F23", X"61", '1'),
      (X"9F23", X"13", '1'),
      (X"9F23", X"61", '1'),
      (X"9F23", X"09", '1'),
      (X"9F23", X"61", '1'),
      (X"9F23", X"03", '1'),
      (X"9F23", X"61", '1'),
      (X"9F23", X"20", '1'),
      (X"9F23", X"61", '1'),
      (X"9F23", X"16", '1'),
      (X"9F23", X"61", '1'),
      (X"9F23", X"32", '1'),
      (X"9F23", X"61", '1'),
      (X"9F23", X"20", '1'),
      (X"9F23", X"61", '1'),
      (X"9F23", X"2A", '1'), -- 0x00150
      (X"9F23", X"61", '1'),
      (X"9F23", X"2A", '1'),
      (X"9F23", X"61", '1'),
      (X"9F23", X"2A", '1'),
      (X"9F23", X"61", '1'),
      (X"9F23", X"2A", '1'),
      (X"9F23", X"61", '1'),

      (X"9F20", X"00", '1'),
      (X"9F21", X"02", '1'), -- Set address to 0x00200
      (X"9F23", X"20", '1'), -- 0x00200
      (X"9F23", X"63", '1'),
      (X"9F23", X"20", '1'),
      (X"9F23", X"63", '1'),
      (X"9F23", X"5F", '1'),
      (X"9F23", X"63", '1'),
      (X"9F23", X"A0", '1'),
      (X"9F23", X"63", '1'),
      (X"9F23", X"A0", '1'),
      (X"9F23", X"63", '1'),
      (X"9F23", X"20", '1'),
      (X"9F23", X"63", '1'),
      (X"9F23", X"A0", '1'),
      (X"9F23", X"63", '1'),
      (X"9F23", X"A0", '1'),
      (X"9F23", X"63", '1'),
      (X"9F23", X"69", '1'), -- 0x00210
      (X"9F23", X"63", '1'),

      (X"9F20", X"00", '1'),
      (X"9F21", X"03", '1'), -- Set address to 0x00300
      (X"9F23", X"20", '1'), -- 0x00300
      (X"9F23", X"65", '1'),
      (X"9F23", X"20", '1'),
      (X"9F23", X"65", '1'),
      (X"9F23", X"20", '1'),
      (X"9F23", X"65", '1'),
      (X"9F23", X"20", '1'),
      (X"9F23", X"65", '1'),
      (X"9F23", X"A0", '1'),
      (X"9F23", X"65", '1'),
      (X"9F23", X"20", '1'),
      (X"9F23", X"65", '1'),
      (X"9F23", X"A0", '1'),
      (X"9F23", X"65", '1'),
      (X"9F23", X"20", '1'),
      (X"9F23", X"61", '1'),
      (X"9F23", X"20", '1'), -- 0x00310
      (X"9F23", X"61", '1'),
      (X"9F23", X"20", '1'),
      (X"9F23", X"61", '1'),
      (X"9F23", X"20", '1'),
      (X"9F23", X"61", '1'),
      (X"9F23", X"20", '1'),
      (X"9F23", X"61", '1'),
      (X"9F23", X"35", '1'),
      (X"9F23", X"61", '1'),
      (X"9F23", X"31", '1'),
      (X"9F23", X"61", '1'),
      (X"9F23", X"32", '1'),
      (X"9F23", X"61", '1'),
      (X"9F23", X"0B", '1'),
      (X"9F23", X"61", '1'),
      (X"9F23", X"20", '1'), -- 0x00320
      (X"9F23", X"61", '1'),
      (X"9F23", X"08", '1'),
      (X"9F23", X"61", '1'),
      (X"9F23", X"09", '1'),
      (X"9F23", X"61", '1'),
      (X"9F23", X"07", '1'),
      (X"9F23", X"61", '1'),
      (X"9F23", X"08", '1'),
      (X"9F23", X"61", '1'),
      (X"9F23", X"20", '1'),
      (X"9F23", X"61", '1'),
      (X"9F23", X"12", '1'),
      (X"9F23", X"61", '1'),
      (X"9F23", X"01", '1'),
      (X"9F23", X"61", '1'),
      (X"9F23", X"0D", '1'), -- 0x00330
      (X"9F23", X"61", '1'),

      (X"9F20", X"00", '1'),
      (X"9F21", X"04", '1'), -- Set address to 0x00400
      (X"9F23", X"20", '1'), -- 0x00400
      (X"9F23", X"67", '1'),
      (X"9F23", X"20", '1'),
      (X"9F23", X"67", '1'),
      (X"9F23", X"E9", '1'),
      (X"9F23", X"67", '1'),
      (X"9F23", X"A0", '1'),
      (X"9F23", X"67", '1'),
      (X"9F23", X"A0", '1'),
      (X"9F23", X"67", '1'),
      (X"9F23", X"20", '1'),
      (X"9F23", X"67", '1'),
      (X"9F23", X"A0", '1'),
      (X"9F23", X"67", '1'),
      (X"9F23", X"A0", '1'),
      (X"9F23", X"67", '1'),
      (X"9F23", X"DF", '1'), -- 0x00410
      (X"9F23", X"67", '1'),

      (X"9F20", X"00", '1'),
      (X"9F21", X"05", '1'), -- Set address to 0x00500
      (X"9F23", X"20", '1'), -- 0x00500
      (X"9F23", X"68", '1'),
      (X"9F23", X"E9", '1'),
      (X"9F23", X"68", '1'),
      (X"9F23", X"A0", '1'),
      (X"9F23", X"68", '1'),
      (X"9F23", X"A0", '1'),
      (X"9F23", X"68", '1'),
      (X"9F23", X"69", '1'),
      (X"9F23", X"68", '1'),
      (X"9F23", X"20", '1'),
      (X"9F23", X"68", '1'),
      (X"9F23", X"5F", '1'),
      (X"9F23", X"68", '1'),
      (X"9F23", X"A0", '1'),
      (X"9F23", X"68", '1'),
      (X"9F23", X"A0", '1'), -- 0x00510
      (X"9F23", X"68", '1'),
      (X"9F23", X"DF", '1'),
      (X"9F23", X"68", '1'),
      (X"9F23", X"20", '1'),
      (X"9F23", X"61", '1'),
      (X"9F23", X"20", '1'),
      (X"9F23", X"61", '1'),
      (X"9F23", X"33", '1'),
      (X"9F23", X"61", '1'),
      (X"9F23", X"38", '1'),
      (X"9F23", X"61", '1'),
      (X"9F23", X"36", '1'),
      (X"9F23", X"61", '1'),
      (X"9F23", X"35", '1'),
      (X"9F23", X"61", '1'),
      (X"9F23", X"35", '1'), -- 0x00520
      (X"9F23", X"61", '1'),
      (X"9F23", X"20", '1'),
      (X"9F23", X"61", '1'),
      (X"9F23", X"02", '1'),
      (X"9F23", X"61", '1'),
      (X"9F23", X"01", '1'),
      (X"9F23", X"61", '1'),
      (X"9F23", X"13", '1'),
      (X"9F23", X"61", '1'),
      (X"9F23", X"09", '1'),
      (X"9F23", X"61", '1'),
      (X"9F23", X"03", '1'),
      (X"9F23", X"61", '1'),
      (X"9F23", X"20", '1'),
      (X"9F23", X"61", '1'),
      (X"9F23", X"02", '1'), -- 0x00530
      (X"9F23", X"61", '1'),
      (X"9F23", X"19", '1'),
      (X"9F23", X"61", '1'),
      (X"9F23", X"14", '1'),
      (X"9F23", X"61", '1'),
      (X"9F23", X"05", '1'),
      (X"9F23", X"61", '1'),
      (X"9F23", X"13", '1'),
      (X"9F23", X"61", '1'),
      (X"9F23", X"20", '1'),
      (X"9F23", X"61", '1'),
      (X"9F23", X"06", '1'),
      (X"9F23", X"61", '1'),
      (X"9F23", X"12", '1'),
      (X"9F23", X"61", '1'),
      (X"9F23", X"05", '1'), -- 0x00540
      (X"9F23", X"61", '1'),
      (X"9F23", X"05", '1'),
      (X"9F23", X"61", '1'),

      (X"9F20", X"00", '1'),
      (X"9F21", X"06", '1'), -- Set address to 0x00600
      (X"9F23", X"E9", '1'), -- 0x00600
      (X"9F23", X"62", '1'),
      (X"9F23", X"A0", '1'),
      (X"9F23", X"62", '1'),
      (X"9F23", X"A0", '1'),
      (X"9F23", X"62", '1'),
      (X"9F23", X"69", '1'),
      (X"9F23", X"62", '1'),
      (X"9F23", X"20", '1'),
      (X"9F23", X"62", '1'),
      (X"9F23", X"20", '1'),
      (X"9F23", X"62", '1'),
      (X"9F23", X"20", '1'),
      (X"9F23", X"62", '1'),
      (X"9F23", X"5F", '1'),
      (X"9F23", X"62", '1'),
      (X"9F23", X"A0", '1'), -- 0x00610
      (X"9F23", X"62", '1'),
      (X"9F23", X"A0", '1'),
      (X"9F23", X"62", '1'),
      (X"9F23", X"DF", '1'),
      (X"9F23", X"62", '1'),

      (X"9F20", X"00", '1'),
      (X"9F21", X"08", '1'), -- Set address to 0x00800
      (X"9F23", X"12", '1'), -- 0x00800
      (X"9F23", X"61", '1'),
      (X"9F23", X"05", '1'),
      (X"9F23", X"61", '1'),
      (X"9F23", X"01", '1'),
      (X"9F23", X"61", '1'),
      (X"9F23", X"04", '1'),
      (X"9F23", X"61", '1'),
      (X"9F23", X"19", '1'),
      (X"9F23", X"61", '1'),
      (X"9F23", X"2E", '1'),
      (X"9F23", X"61", '1'),

      -- The second part is the tile map, i.e. the font
      (X"9F20", X"00", '1'),
      (X"9F21", X"F8", '1'), -- Set address to 0x0F800
      (X"9F23", X"3C", '1'), -- 0x0F800
      (X"9F23", X"66", '1'),
      (X"9F23", X"6E", '1'),
      (X"9F23", X"6E", '1'),
      (X"9F23", X"60", '1'),
      (X"9F23", X"62", '1'),
      (X"9F23", X"3C", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"18", '1'),
      (X"9F23", X"3C", '1'),
      (X"9F23", X"66", '1'),
      (X"9F23", X"7E", '1'),
      (X"9F23", X"66", '1'),
      (X"9F23", X"66", '1'),
      (X"9F23", X"66", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"7C", '1'),
      (X"9F23", X"66", '1'),
      (X"9F23", X"66", '1'),
      (X"9F23", X"7C", '1'),
      (X"9F23", X"66", '1'),
      (X"9F23", X"66", '1'),
      (X"9F23", X"7C", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"3C", '1'),
      (X"9F23", X"66", '1'),
      (X"9F23", X"60", '1'),
      (X"9F23", X"60", '1'),
      (X"9F23", X"60", '1'),
      (X"9F23", X"66", '1'),
      (X"9F23", X"3C", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"78", '1'),
      (X"9F23", X"6C", '1'),
      (X"9F23", X"66", '1'),
      (X"9F23", X"66", '1'),
      (X"9F23", X"66", '1'),
      (X"9F23", X"6C", '1'),
      (X"9F23", X"78", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"7E", '1'),
      (X"9F23", X"60", '1'),
      (X"9F23", X"60", '1'),
      (X"9F23", X"78", '1'),
      (X"9F23", X"60", '1'),
      (X"9F23", X"60", '1'),
      (X"9F23", X"7E", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"7E", '1'),
      (X"9F23", X"60", '1'),
      (X"9F23", X"60", '1'),
      (X"9F23", X"78", '1'),
      (X"9F23", X"60", '1'),
      (X"9F23", X"60", '1'),
      (X"9F23", X"60", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"3C", '1'),
      (X"9F23", X"66", '1'),
      (X"9F23", X"60", '1'),
      (X"9F23", X"6E", '1'),
      (X"9F23", X"66", '1'),
      (X"9F23", X"66", '1'),
      (X"9F23", X"3C", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"66", '1'),
      (X"9F23", X"66", '1'),
      (X"9F23", X"66", '1'),
      (X"9F23", X"7E", '1'),
      (X"9F23", X"66", '1'),
      (X"9F23", X"66", '1'),
      (X"9F23", X"66", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"3C", '1'),
      (X"9F23", X"18", '1'),
      (X"9F23", X"18", '1'),
      (X"9F23", X"18", '1'),
      (X"9F23", X"18", '1'),
      (X"9F23", X"18", '1'),
      (X"9F23", X"3C", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"1E", '1'),
      (X"9F23", X"0C", '1'),
      (X"9F23", X"0C", '1'),
      (X"9F23", X"0C", '1'),
      (X"9F23", X"0C", '1'),
      (X"9F23", X"6C", '1'),
      (X"9F23", X"38", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"66", '1'),
      (X"9F23", X"6C", '1'),
      (X"9F23", X"78", '1'),
      (X"9F23", X"70", '1'),
      (X"9F23", X"78", '1'),
      (X"9F23", X"6C", '1'),
      (X"9F23", X"66", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"60", '1'),
      (X"9F23", X"60", '1'),
      (X"9F23", X"60", '1'),
      (X"9F23", X"60", '1'),
      (X"9F23", X"60", '1'),
      (X"9F23", X"60", '1'),
      (X"9F23", X"7E", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"63", '1'),
      (X"9F23", X"77", '1'),
      (X"9F23", X"7F", '1'),
      (X"9F23", X"6B", '1'),
      (X"9F23", X"63", '1'),
      (X"9F23", X"63", '1'),
      (X"9F23", X"63", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"66", '1'),
      (X"9F23", X"76", '1'),
      (X"9F23", X"7E", '1'),
      (X"9F23", X"7E", '1'),
      (X"9F23", X"6E", '1'),
      (X"9F23", X"66", '1'),
      (X"9F23", X"66", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"3C", '1'),
      (X"9F23", X"66", '1'),
      (X"9F23", X"66", '1'),
      (X"9F23", X"66", '1'),
      (X"9F23", X"66", '1'),
      (X"9F23", X"66", '1'),
      (X"9F23", X"3C", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"7C", '1'),
      (X"9F23", X"66", '1'),
      (X"9F23", X"66", '1'),
      (X"9F23", X"7C", '1'),
      (X"9F23", X"60", '1'),
      (X"9F23", X"60", '1'),
      (X"9F23", X"60", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"3C", '1'),
      (X"9F23", X"66", '1'),
      (X"9F23", X"66", '1'),
      (X"9F23", X"66", '1'),
      (X"9F23", X"66", '1'),
      (X"9F23", X"3C", '1'),
      (X"9F23", X"0E", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"7C", '1'),
      (X"9F23", X"66", '1'),
      (X"9F23", X"66", '1'),
      (X"9F23", X"7C", '1'),
      (X"9F23", X"78", '1'),
      (X"9F23", X"6C", '1'),
      (X"9F23", X"66", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"3C", '1'),
      (X"9F23", X"66", '1'),
      (X"9F23", X"60", '1'),
      (X"9F23", X"3C", '1'),
      (X"9F23", X"06", '1'),
      (X"9F23", X"66", '1'),
      (X"9F23", X"3C", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"7E", '1'),
      (X"9F23", X"18", '1'),
      (X"9F23", X"18", '1'),
      (X"9F23", X"18", '1'),
      (X"9F23", X"18", '1'),
      (X"9F23", X"18", '1'),
      (X"9F23", X"18", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"66", '1'),
      (X"9F23", X"66", '1'),
      (X"9F23", X"66", '1'),
      (X"9F23", X"66", '1'),
      (X"9F23", X"66", '1'),
      (X"9F23", X"66", '1'),
      (X"9F23", X"3C", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"66", '1'),
      (X"9F23", X"66", '1'),
      (X"9F23", X"66", '1'),
      (X"9F23", X"66", '1'),
      (X"9F23", X"66", '1'),
      (X"9F23", X"3C", '1'),
      (X"9F23", X"18", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"63", '1'),
      (X"9F23", X"63", '1'),
      (X"9F23", X"63", '1'),
      (X"9F23", X"6B", '1'),
      (X"9F23", X"7F", '1'),
      (X"9F23", X"77", '1'),
      (X"9F23", X"63", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"66", '1'),
      (X"9F23", X"66", '1'),
      (X"9F23", X"3C", '1'),
      (X"9F23", X"18", '1'),
      (X"9F23", X"3C", '1'),
      (X"9F23", X"66", '1'),
      (X"9F23", X"66", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"66", '1'),
      (X"9F23", X"66", '1'),
      (X"9F23", X"66", '1'),
      (X"9F23", X"3C", '1'),
      (X"9F23", X"18", '1'),
      (X"9F23", X"18", '1'),
      (X"9F23", X"18", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"7E", '1'),
      (X"9F23", X"06", '1'),
      (X"9F23", X"0C", '1'),
      (X"9F23", X"18", '1'),
      (X"9F23", X"30", '1'),
      (X"9F23", X"60", '1'),
      (X"9F23", X"7E", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"3C", '1'),
      (X"9F23", X"30", '1'),
      (X"9F23", X"30", '1'),
      (X"9F23", X"30", '1'),
      (X"9F23", X"30", '1'),
      (X"9F23", X"30", '1'),
      (X"9F23", X"3C", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"0C", '1'),
      (X"9F23", X"12", '1'),
      (X"9F23", X"30", '1'),
      (X"9F23", X"7C", '1'),
      (X"9F23", X"30", '1'),
      (X"9F23", X"62", '1'),
      (X"9F23", X"FC", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"3C", '1'),
      (X"9F23", X"0C", '1'),
      (X"9F23", X"0C", '1'),
      (X"9F23", X"0C", '1'),
      (X"9F23", X"0C", '1'),
      (X"9F23", X"0C", '1'),
      (X"9F23", X"3C", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"18", '1'),
      (X"9F23", X"3C", '1'),
      (X"9F23", X"7E", '1'),
      (X"9F23", X"18", '1'),
      (X"9F23", X"18", '1'),
      (X"9F23", X"18", '1'),
      (X"9F23", X"18", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"10", '1'),
      (X"9F23", X"30", '1'),
      (X"9F23", X"7F", '1'),
      (X"9F23", X"7F", '1'),
      (X"9F23", X"30", '1'),
      (X"9F23", X"10", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'), -- 0x0F900
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"18", '1'),
      (X"9F23", X"18", '1'),
      (X"9F23", X"18", '1'),
      (X"9F23", X"18", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"18", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"66", '1'),
      (X"9F23", X"66", '1'),
      (X"9F23", X"66", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"66", '1'),
      (X"9F23", X"66", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"66", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"66", '1'),
      (X"9F23", X"66", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"18", '1'),
      (X"9F23", X"3E", '1'),
      (X"9F23", X"60", '1'),
      (X"9F23", X"3C", '1'),
      (X"9F23", X"06", '1'),
      (X"9F23", X"7C", '1'),
      (X"9F23", X"18", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"62", '1'),
      (X"9F23", X"66", '1'),
      (X"9F23", X"0C", '1'),
      (X"9F23", X"18", '1'),
      (X"9F23", X"30", '1'),
      (X"9F23", X"66", '1'),
      (X"9F23", X"46", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"3C", '1'),
      (X"9F23", X"66", '1'),
      (X"9F23", X"3C", '1'),
      (X"9F23", X"38", '1'),
      (X"9F23", X"67", '1'),
      (X"9F23", X"66", '1'),
      (X"9F23", X"3F", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"06", '1'),
      (X"9F23", X"0C", '1'),
      (X"9F23", X"18", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"0C", '1'),
      (X"9F23", X"18", '1'),
      (X"9F23", X"30", '1'),
      (X"9F23", X"30", '1'),
      (X"9F23", X"30", '1'),
      (X"9F23", X"18", '1'),
      (X"9F23", X"0C", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"30", '1'),
      (X"9F23", X"18", '1'),
      (X"9F23", X"0C", '1'),
      (X"9F23", X"0C", '1'),
      (X"9F23", X"0C", '1'),
      (X"9F23", X"18", '1'),
      (X"9F23", X"30", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"66", '1'),
      (X"9F23", X"3C", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"3C", '1'),
      (X"9F23", X"66", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"18", '1'),
      (X"9F23", X"18", '1'),
      (X"9F23", X"7E", '1'),
      (X"9F23", X"18", '1'),
      (X"9F23", X"18", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"18", '1'),
      (X"9F23", X"18", '1'),
      (X"9F23", X"30", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"7E", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"18", '1'),
      (X"9F23", X"18", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"03", '1'),
      (X"9F23", X"06", '1'),
      (X"9F23", X"0C", '1'),
      (X"9F23", X"18", '1'),
      (X"9F23", X"30", '1'),
      (X"9F23", X"60", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"3C", '1'),
      (X"9F23", X"66", '1'),
      (X"9F23", X"6E", '1'),
      (X"9F23", X"76", '1'),
      (X"9F23", X"66", '1'),
      (X"9F23", X"66", '1'),
      (X"9F23", X"3C", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"18", '1'),
      (X"9F23", X"18", '1'),
      (X"9F23", X"38", '1'),
      (X"9F23", X"18", '1'),
      (X"9F23", X"18", '1'),
      (X"9F23", X"18", '1'),
      (X"9F23", X"7E", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"3C", '1'),
      (X"9F23", X"66", '1'),
      (X"9F23", X"06", '1'),
      (X"9F23", X"0C", '1'),
      (X"9F23", X"30", '1'),
      (X"9F23", X"60", '1'),
      (X"9F23", X"7E", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"3C", '1'),
      (X"9F23", X"66", '1'),
      (X"9F23", X"06", '1'),
      (X"9F23", X"1C", '1'),
      (X"9F23", X"06", '1'),
      (X"9F23", X"66", '1'),
      (X"9F23", X"3C", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"06", '1'),
      (X"9F23", X"0E", '1'),
      (X"9F23", X"1E", '1'),
      (X"9F23", X"66", '1'),
      (X"9F23", X"7F", '1'),
      (X"9F23", X"06", '1'),
      (X"9F23", X"06", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"7E", '1'),
      (X"9F23", X"60", '1'),
      (X"9F23", X"7C", '1'),
      (X"9F23", X"06", '1'),
      (X"9F23", X"06", '1'),
      (X"9F23", X"66", '1'),
      (X"9F23", X"3C", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"3C", '1'),
      (X"9F23", X"66", '1'),
      (X"9F23", X"60", '1'),
      (X"9F23", X"7C", '1'),
      (X"9F23", X"66", '1'),
      (X"9F23", X"66", '1'),
      (X"9F23", X"3C", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"7E", '1'),
      (X"9F23", X"66", '1'),
      (X"9F23", X"0C", '1'),
      (X"9F23", X"18", '1'),
      (X"9F23", X"18", '1'),
      (X"9F23", X"18", '1'),
      (X"9F23", X"18", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"3C", '1'),
      (X"9F23", X"66", '1'),
      (X"9F23", X"66", '1'),
      (X"9F23", X"3C", '1'),
      (X"9F23", X"66", '1'),
      (X"9F23", X"66", '1'),
      (X"9F23", X"3C", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"3C", '1'),
      (X"9F23", X"66", '1'),
      (X"9F23", X"66", '1'),
      (X"9F23", X"3E", '1'),
      (X"9F23", X"06", '1'),
      (X"9F23", X"66", '1'),
      (X"9F23", X"3C", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"18", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"18", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"18", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"18", '1'),
      (X"9F23", X"18", '1'),
      (X"9F23", X"30", '1'),
      (X"9F23", X"0E", '1'),
      (X"9F23", X"18", '1'),
      (X"9F23", X"30", '1'),
      (X"9F23", X"60", '1'),
      (X"9F23", X"30", '1'),
      (X"9F23", X"18", '1'),
      (X"9F23", X"0E", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"7E", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"7E", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"70", '1'),
      (X"9F23", X"18", '1'),
      (X"9F23", X"0C", '1'),
      (X"9F23", X"06", '1'),
      (X"9F23", X"0C", '1'),
      (X"9F23", X"18", '1'),
      (X"9F23", X"70", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"3C", '1'),
      (X"9F23", X"66", '1'),
      (X"9F23", X"06", '1'),
      (X"9F23", X"0C", '1'),
      (X"9F23", X"18", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"18", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'), -- 0x0FA00
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"08", '1'),
      (X"9F23", X"1C", '1'),
      (X"9F23", X"3E", '1'),
      (X"9F23", X"7F", '1'),
      (X"9F23", X"7F", '1'),
      (X"9F23", X"1C", '1'),
      (X"9F23", X"3E", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"18", '1'),
      (X"9F23", X"18", '1'),
      (X"9F23", X"18", '1'),
      (X"9F23", X"18", '1'),
      (X"9F23", X"18", '1'),
      (X"9F23", X"18", '1'),
      (X"9F23", X"18", '1'),
      (X"9F23", X"18", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"30", '1'),
      (X"9F23", X"30", '1'),
      (X"9F23", X"30", '1'),
      (X"9F23", X"30", '1'),
      (X"9F23", X"30", '1'),
      (X"9F23", X"30", '1'),
      (X"9F23", X"30", '1'),
      (X"9F23", X"30", '1'),
      (X"9F23", X"0C", '1'),
      (X"9F23", X"0C", '1'),
      (X"9F23", X"0C", '1'),
      (X"9F23", X"0C", '1'),
      (X"9F23", X"0C", '1'),
      (X"9F23", X"0C", '1'),
      (X"9F23", X"0C", '1'),
      (X"9F23", X"0C", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"E0", '1'),
      (X"9F23", X"F0", '1'),
      (X"9F23", X"38", '1'),
      (X"9F23", X"18", '1'),
      (X"9F23", X"18", '1'),
      (X"9F23", X"18", '1'),
      (X"9F23", X"18", '1'),
      (X"9F23", X"1C", '1'),
      (X"9F23", X"0F", '1'),
      (X"9F23", X"07", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"18", '1'),
      (X"9F23", X"18", '1'),
      (X"9F23", X"38", '1'),
      (X"9F23", X"F0", '1'),
      (X"9F23", X"E0", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"C0", '1'),
      (X"9F23", X"C0", '1'),
      (X"9F23", X"C0", '1'),
      (X"9F23", X"C0", '1'),
      (X"9F23", X"C0", '1'),
      (X"9F23", X"C0", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"C0", '1'),
      (X"9F23", X"E0", '1'),
      (X"9F23", X"70", '1'),
      (X"9F23", X"38", '1'),
      (X"9F23", X"1C", '1'),
      (X"9F23", X"0E", '1'),
      (X"9F23", X"07", '1'),
      (X"9F23", X"03", '1'),
      (X"9F23", X"03", '1'),
      (X"9F23", X"07", '1'),
      (X"9F23", X"0E", '1'),
      (X"9F23", X"1C", '1'),
      (X"9F23", X"38", '1'),
      (X"9F23", X"70", '1'),
      (X"9F23", X"E0", '1'),
      (X"9F23", X"C0", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"C0", '1'),
      (X"9F23", X"C0", '1'),
      (X"9F23", X"C0", '1'),
      (X"9F23", X"C0", '1'),
      (X"9F23", X"C0", '1'),
      (X"9F23", X"C0", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"03", '1'),
      (X"9F23", X"03", '1'),
      (X"9F23", X"03", '1'),
      (X"9F23", X"03", '1'),
      (X"9F23", X"03", '1'),
      (X"9F23", X"03", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"3C", '1'),
      (X"9F23", X"7E", '1'),
      (X"9F23", X"7E", '1'),
      (X"9F23", X"7E", '1'),
      (X"9F23", X"7E", '1'),
      (X"9F23", X"3C", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"36", '1'),
      (X"9F23", X"7F", '1'),
      (X"9F23", X"7F", '1'),
      (X"9F23", X"7F", '1'),
      (X"9F23", X"3E", '1'),
      (X"9F23", X"1C", '1'),
      (X"9F23", X"08", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"60", '1'),
      (X"9F23", X"60", '1'),
      (X"9F23", X"60", '1'),
      (X"9F23", X"60", '1'),
      (X"9F23", X"60", '1'),
      (X"9F23", X"60", '1'),
      (X"9F23", X"60", '1'),
      (X"9F23", X"60", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"07", '1'),
      (X"9F23", X"0F", '1'),
      (X"9F23", X"1C", '1'),
      (X"9F23", X"18", '1'),
      (X"9F23", X"18", '1'),
      (X"9F23", X"C3", '1'),
      (X"9F23", X"E7", '1'),
      (X"9F23", X"7E", '1'),
      (X"9F23", X"3C", '1'),
      (X"9F23", X"3C", '1'),
      (X"9F23", X"7E", '1'),
      (X"9F23", X"E7", '1'),
      (X"9F23", X"C3", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"3C", '1'),
      (X"9F23", X"7E", '1'),
      (X"9F23", X"66", '1'),
      (X"9F23", X"66", '1'),
      (X"9F23", X"7E", '1'),
      (X"9F23", X"3C", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"18", '1'),
      (X"9F23", X"18", '1'),
      (X"9F23", X"66", '1'),
      (X"9F23", X"66", '1'),
      (X"9F23", X"18", '1'),
      (X"9F23", X"18", '1'),
      (X"9F23", X"3C", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"06", '1'),
      (X"9F23", X"06", '1'),
      (X"9F23", X"06", '1'),
      (X"9F23", X"06", '1'),
      (X"9F23", X"06", '1'),
      (X"9F23", X"06", '1'),
      (X"9F23", X"06", '1'),
      (X"9F23", X"06", '1'),
      (X"9F23", X"08", '1'),
      (X"9F23", X"1C", '1'),
      (X"9F23", X"3E", '1'),
      (X"9F23", X"7F", '1'),
      (X"9F23", X"3E", '1'),
      (X"9F23", X"1C", '1'),
      (X"9F23", X"08", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"18", '1'),
      (X"9F23", X"18", '1'),
      (X"9F23", X"18", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"18", '1'),
      (X"9F23", X"18", '1'),
      (X"9F23", X"18", '1'),
      (X"9F23", X"C0", '1'),
      (X"9F23", X"C0", '1'),
      (X"9F23", X"30", '1'),
      (X"9F23", X"30", '1'),
      (X"9F23", X"C0", '1'),
      (X"9F23", X"C0", '1'),
      (X"9F23", X"30", '1'),
      (X"9F23", X"30", '1'),
      (X"9F23", X"18", '1'),
      (X"9F23", X"18", '1'),
      (X"9F23", X"18", '1'),
      (X"9F23", X"18", '1'),
      (X"9F23", X"18", '1'),
      (X"9F23", X"18", '1'),
      (X"9F23", X"18", '1'),
      (X"9F23", X"18", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"03", '1'),
      (X"9F23", X"3E", '1'),
      (X"9F23", X"76", '1'),
      (X"9F23", X"36", '1'),
      (X"9F23", X"36", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"7F", '1'),
      (X"9F23", X"3F", '1'),
      (X"9F23", X"1F", '1'),
      (X"9F23", X"0F", '1'),
      (X"9F23", X"07", '1'),
      (X"9F23", X"03", '1'),
      (X"9F23", X"01", '1'),
      (X"9F23", X"00", '1'), -- 0x0FB00
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"F0", '1'),
      (X"9F23", X"F0", '1'),
      (X"9F23", X"F0", '1'),
      (X"9F23", X"F0", '1'),
      (X"9F23", X"F0", '1'),
      (X"9F23", X"F0", '1'),
      (X"9F23", X"F0", '1'),
      (X"9F23", X"F0", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"C0", '1'),
      (X"9F23", X"C0", '1'),
      (X"9F23", X"C0", '1'),
      (X"9F23", X"C0", '1'),
      (X"9F23", X"C0", '1'),
      (X"9F23", X"C0", '1'),
      (X"9F23", X"C0", '1'),
      (X"9F23", X"C0", '1'),
      (X"9F23", X"CC", '1'),
      (X"9F23", X"CC", '1'),
      (X"9F23", X"33", '1'),
      (X"9F23", X"33", '1'),
      (X"9F23", X"CC", '1'),
      (X"9F23", X"CC", '1'),
      (X"9F23", X"33", '1'),
      (X"9F23", X"33", '1'),
      (X"9F23", X"03", '1'),
      (X"9F23", X"03", '1'),
      (X"9F23", X"03", '1'),
      (X"9F23", X"03", '1'),
      (X"9F23", X"03", '1'),
      (X"9F23", X"03", '1'),
      (X"9F23", X"03", '1'),
      (X"9F23", X"03", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"CC", '1'),
      (X"9F23", X"CC", '1'),
      (X"9F23", X"33", '1'),
      (X"9F23", X"33", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FE", '1'),
      (X"9F23", X"FC", '1'),
      (X"9F23", X"F8", '1'),
      (X"9F23", X"F0", '1'),
      (X"9F23", X"E0", '1'),
      (X"9F23", X"C0", '1'),
      (X"9F23", X"80", '1'),
      (X"9F23", X"03", '1'),
      (X"9F23", X"03", '1'),
      (X"9F23", X"03", '1'),
      (X"9F23", X"03", '1'),
      (X"9F23", X"03", '1'),
      (X"9F23", X"03", '1'),
      (X"9F23", X"03", '1'),
      (X"9F23", X"03", '1'),
      (X"9F23", X"18", '1'),
      (X"9F23", X"18", '1'),
      (X"9F23", X"18", '1'),
      (X"9F23", X"1F", '1'),
      (X"9F23", X"1F", '1'),
      (X"9F23", X"18", '1'),
      (X"9F23", X"18", '1'),
      (X"9F23", X"18", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"0F", '1'),
      (X"9F23", X"0F", '1'),
      (X"9F23", X"0F", '1'),
      (X"9F23", X"0F", '1'),
      (X"9F23", X"18", '1'),
      (X"9F23", X"18", '1'),
      (X"9F23", X"18", '1'),
      (X"9F23", X"1F", '1'),
      (X"9F23", X"1F", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"F8", '1'),
      (X"9F23", X"F8", '1'),
      (X"9F23", X"18", '1'),
      (X"9F23", X"18", '1'),
      (X"9F23", X"18", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"1F", '1'),
      (X"9F23", X"1F", '1'),
      (X"9F23", X"18", '1'),
      (X"9F23", X"18", '1'),
      (X"9F23", X"18", '1'),
      (X"9F23", X"18", '1'),
      (X"9F23", X"18", '1'),
      (X"9F23", X"18", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"18", '1'),
      (X"9F23", X"18", '1'),
      (X"9F23", X"18", '1'),
      (X"9F23", X"18", '1'),
      (X"9F23", X"18", '1'),
      (X"9F23", X"18", '1'),
      (X"9F23", X"F8", '1'),
      (X"9F23", X"F8", '1'),
      (X"9F23", X"18", '1'),
      (X"9F23", X"18", '1'),
      (X"9F23", X"18", '1'),
      (X"9F23", X"C0", '1'),
      (X"9F23", X"C0", '1'),
      (X"9F23", X"C0", '1'),
      (X"9F23", X"C0", '1'),
      (X"9F23", X"C0", '1'),
      (X"9F23", X"C0", '1'),
      (X"9F23", X"C0", '1'),
      (X"9F23", X"C0", '1'),
      (X"9F23", X"E0", '1'),
      (X"9F23", X"E0", '1'),
      (X"9F23", X"E0", '1'),
      (X"9F23", X"E0", '1'),
      (X"9F23", X"E0", '1'),
      (X"9F23", X"E0", '1'),
      (X"9F23", X"E0", '1'),
      (X"9F23", X"E0", '1'),
      (X"9F23", X"07", '1'),
      (X"9F23", X"07", '1'),
      (X"9F23", X"07", '1'),
      (X"9F23", X"07", '1'),
      (X"9F23", X"07", '1'),
      (X"9F23", X"07", '1'),
      (X"9F23", X"07", '1'),
      (X"9F23", X"07", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"03", '1'),
      (X"9F23", X"03", '1'),
      (X"9F23", X"03", '1'),
      (X"9F23", X"03", '1'),
      (X"9F23", X"03", '1'),
      (X"9F23", X"03", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"F0", '1'),
      (X"9F23", X"F0", '1'),
      (X"9F23", X"F0", '1'),
      (X"9F23", X"F0", '1'),
      (X"9F23", X"0F", '1'),
      (X"9F23", X"0F", '1'),
      (X"9F23", X"0F", '1'),
      (X"9F23", X"0F", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"18", '1'),
      (X"9F23", X"18", '1'),
      (X"9F23", X"18", '1'),
      (X"9F23", X"F8", '1'),
      (X"9F23", X"F8", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"F0", '1'),
      (X"9F23", X"F0", '1'),
      (X"9F23", X"F0", '1'),
      (X"9F23", X"F0", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"F0", '1'),
      (X"9F23", X"F0", '1'),
      (X"9F23", X"F0", '1'),
      (X"9F23", X"F0", '1'),
      (X"9F23", X"0F", '1'),
      (X"9F23", X"0F", '1'),
      (X"9F23", X"0F", '1'),
      (X"9F23", X"0F", '1'),
      (X"9F23", X"C3", '1'), -- 0x0FC00
      (X"9F23", X"99", '1'),
      (X"9F23", X"91", '1'),
      (X"9F23", X"91", '1'),
      (X"9F23", X"9F", '1'),
      (X"9F23", X"9D", '1'),
      (X"9F23", X"C3", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"E7", '1'),
      (X"9F23", X"C3", '1'),
      (X"9F23", X"99", '1'),
      (X"9F23", X"81", '1'),
      (X"9F23", X"99", '1'),
      (X"9F23", X"99", '1'),
      (X"9F23", X"99", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"83", '1'),
      (X"9F23", X"99", '1'),
      (X"9F23", X"99", '1'),
      (X"9F23", X"83", '1'),
      (X"9F23", X"99", '1'),
      (X"9F23", X"99", '1'),
      (X"9F23", X"83", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"C3", '1'),
      (X"9F23", X"99", '1'),
      (X"9F23", X"9F", '1'),
      (X"9F23", X"9F", '1'),
      (X"9F23", X"9F", '1'),
      (X"9F23", X"99", '1'),
      (X"9F23", X"C3", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"87", '1'),
      (X"9F23", X"93", '1'),
      (X"9F23", X"99", '1'),
      (X"9F23", X"99", '1'),
      (X"9F23", X"99", '1'),
      (X"9F23", X"93", '1'),
      (X"9F23", X"87", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"81", '1'),
      (X"9F23", X"9F", '1'),
      (X"9F23", X"9F", '1'),
      (X"9F23", X"87", '1'),
      (X"9F23", X"9F", '1'),
      (X"9F23", X"9F", '1'),
      (X"9F23", X"81", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"81", '1'),
      (X"9F23", X"9F", '1'),
      (X"9F23", X"9F", '1'),
      (X"9F23", X"87", '1'),
      (X"9F23", X"9F", '1'),
      (X"9F23", X"9F", '1'),
      (X"9F23", X"9F", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"C3", '1'),
      (X"9F23", X"99", '1'),
      (X"9F23", X"9F", '1'),
      (X"9F23", X"91", '1'),
      (X"9F23", X"99", '1'),
      (X"9F23", X"99", '1'),
      (X"9F23", X"C3", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"99", '1'),
      (X"9F23", X"99", '1'),
      (X"9F23", X"99", '1'),
      (X"9F23", X"81", '1'),
      (X"9F23", X"99", '1'),
      (X"9F23", X"99", '1'),
      (X"9F23", X"99", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"C3", '1'),
      (X"9F23", X"E7", '1'),
      (X"9F23", X"E7", '1'),
      (X"9F23", X"E7", '1'),
      (X"9F23", X"E7", '1'),
      (X"9F23", X"E7", '1'),
      (X"9F23", X"C3", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"E1", '1'),
      (X"9F23", X"F3", '1'),
      (X"9F23", X"F3", '1'),
      (X"9F23", X"F3", '1'),
      (X"9F23", X"F3", '1'),
      (X"9F23", X"93", '1'),
      (X"9F23", X"C7", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"99", '1'),
      (X"9F23", X"93", '1'),
      (X"9F23", X"87", '1'),
      (X"9F23", X"8F", '1'),
      (X"9F23", X"87", '1'),
      (X"9F23", X"93", '1'),
      (X"9F23", X"99", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"9F", '1'),
      (X"9F23", X"9F", '1'),
      (X"9F23", X"9F", '1'),
      (X"9F23", X"9F", '1'),
      (X"9F23", X"9F", '1'),
      (X"9F23", X"9F", '1'),
      (X"9F23", X"81", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"9C", '1'),
      (X"9F23", X"88", '1'),
      (X"9F23", X"80", '1'),
      (X"9F23", X"94", '1'),
      (X"9F23", X"9C", '1'),
      (X"9F23", X"9C", '1'),
      (X"9F23", X"9C", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"99", '1'),
      (X"9F23", X"89", '1'),
      (X"9F23", X"81", '1'),
      (X"9F23", X"81", '1'),
      (X"9F23", X"91", '1'),
      (X"9F23", X"99", '1'),
      (X"9F23", X"99", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"C3", '1'),
      (X"9F23", X"99", '1'),
      (X"9F23", X"99", '1'),
      (X"9F23", X"99", '1'),
      (X"9F23", X"99", '1'),
      (X"9F23", X"99", '1'),
      (X"9F23", X"C3", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"83", '1'),
      (X"9F23", X"99", '1'),
      (X"9F23", X"99", '1'),
      (X"9F23", X"83", '1'),
      (X"9F23", X"9F", '1'),
      (X"9F23", X"9F", '1'),
      (X"9F23", X"9F", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"C3", '1'),
      (X"9F23", X"99", '1'),
      (X"9F23", X"99", '1'),
      (X"9F23", X"99", '1'),
      (X"9F23", X"99", '1'),
      (X"9F23", X"C3", '1'),
      (X"9F23", X"F1", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"83", '1'),
      (X"9F23", X"99", '1'),
      (X"9F23", X"99", '1'),
      (X"9F23", X"83", '1'),
      (X"9F23", X"87", '1'),
      (X"9F23", X"93", '1'),
      (X"9F23", X"99", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"C3", '1'),
      (X"9F23", X"99", '1'),
      (X"9F23", X"9F", '1'),
      (X"9F23", X"C3", '1'),
      (X"9F23", X"F9", '1'),
      (X"9F23", X"99", '1'),
      (X"9F23", X"C3", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"81", '1'),
      (X"9F23", X"E7", '1'),
      (X"9F23", X"E7", '1'),
      (X"9F23", X"E7", '1'),
      (X"9F23", X"E7", '1'),
      (X"9F23", X"E7", '1'),
      (X"9F23", X"E7", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"99", '1'),
      (X"9F23", X"99", '1'),
      (X"9F23", X"99", '1'),
      (X"9F23", X"99", '1'),
      (X"9F23", X"99", '1'),
      (X"9F23", X"99", '1'),
      (X"9F23", X"C3", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"99", '1'),
      (X"9F23", X"99", '1'),
      (X"9F23", X"99", '1'),
      (X"9F23", X"99", '1'),
      (X"9F23", X"99", '1'),
      (X"9F23", X"C3", '1'),
      (X"9F23", X"E7", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"9C", '1'),
      (X"9F23", X"9C", '1'),
      (X"9F23", X"9C", '1'),
      (X"9F23", X"94", '1'),
      (X"9F23", X"80", '1'),
      (X"9F23", X"88", '1'),
      (X"9F23", X"9C", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"99", '1'),
      (X"9F23", X"99", '1'),
      (X"9F23", X"C3", '1'),
      (X"9F23", X"E7", '1'),
      (X"9F23", X"C3", '1'),
      (X"9F23", X"99", '1'),
      (X"9F23", X"99", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"99", '1'),
      (X"9F23", X"99", '1'),
      (X"9F23", X"99", '1'),
      (X"9F23", X"C3", '1'),
      (X"9F23", X"E7", '1'),
      (X"9F23", X"E7", '1'),
      (X"9F23", X"E7", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"81", '1'),
      (X"9F23", X"F9", '1'),
      (X"9F23", X"F3", '1'),
      (X"9F23", X"E7", '1'),
      (X"9F23", X"CF", '1'),
      (X"9F23", X"9F", '1'),
      (X"9F23", X"81", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"C3", '1'),
      (X"9F23", X"CF", '1'),
      (X"9F23", X"CF", '1'),
      (X"9F23", X"CF", '1'),
      (X"9F23", X"CF", '1'),
      (X"9F23", X"CF", '1'),
      (X"9F23", X"C3", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"F3", '1'),
      (X"9F23", X"ED", '1'),
      (X"9F23", X"CF", '1'),
      (X"9F23", X"83", '1'),
      (X"9F23", X"CF", '1'),
      (X"9F23", X"9D", '1'),
      (X"9F23", X"03", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"C3", '1'),
      (X"9F23", X"F3", '1'),
      (X"9F23", X"F3", '1'),
      (X"9F23", X"F3", '1'),
      (X"9F23", X"F3", '1'),
      (X"9F23", X"F3", '1'),
      (X"9F23", X"C3", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"E7", '1'),
      (X"9F23", X"C3", '1'),
      (X"9F23", X"81", '1'),
      (X"9F23", X"E7", '1'),
      (X"9F23", X"E7", '1'),
      (X"9F23", X"E7", '1'),
      (X"9F23", X"E7", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"EF", '1'),
      (X"9F23", X"CF", '1'),
      (X"9F23", X"80", '1'),
      (X"9F23", X"80", '1'),
      (X"9F23", X"CF", '1'),
      (X"9F23", X"EF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'), -- 0x0FD00
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"E7", '1'),
      (X"9F23", X"E7", '1'),
      (X"9F23", X"E7", '1'),
      (X"9F23", X"E7", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"E7", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"99", '1'),
      (X"9F23", X"99", '1'),
      (X"9F23", X"99", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"99", '1'),
      (X"9F23", X"99", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"99", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"99", '1'),
      (X"9F23", X"99", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"E7", '1'),
      (X"9F23", X"C1", '1'),
      (X"9F23", X"9F", '1'),
      (X"9F23", X"C3", '1'),
      (X"9F23", X"F9", '1'),
      (X"9F23", X"83", '1'),
      (X"9F23", X"E7", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"9D", '1'),
      (X"9F23", X"99", '1'),
      (X"9F23", X"F3", '1'),
      (X"9F23", X"E7", '1'),
      (X"9F23", X"CF", '1'),
      (X"9F23", X"99", '1'),
      (X"9F23", X"B9", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"C3", '1'),
      (X"9F23", X"99", '1'),
      (X"9F23", X"C3", '1'),
      (X"9F23", X"C7", '1'),
      (X"9F23", X"98", '1'),
      (X"9F23", X"99", '1'),
      (X"9F23", X"C0", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"F9", '1'),
      (X"9F23", X"F3", '1'),
      (X"9F23", X"E7", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"F3", '1'),
      (X"9F23", X"E7", '1'),
      (X"9F23", X"CF", '1'),
      (X"9F23", X"CF", '1'),
      (X"9F23", X"CF", '1'),
      (X"9F23", X"E7", '1'),
      (X"9F23", X"F3", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"CF", '1'),
      (X"9F23", X"E7", '1'),
      (X"9F23", X"F3", '1'),
      (X"9F23", X"F3", '1'),
      (X"9F23", X"F3", '1'),
      (X"9F23", X"E7", '1'),
      (X"9F23", X"CF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"99", '1'),
      (X"9F23", X"C3", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"C3", '1'),
      (X"9F23", X"99", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"E7", '1'),
      (X"9F23", X"E7", '1'),
      (X"9F23", X"81", '1'),
      (X"9F23", X"E7", '1'),
      (X"9F23", X"E7", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"E7", '1'),
      (X"9F23", X"E7", '1'),
      (X"9F23", X"CF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"81", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"E7", '1'),
      (X"9F23", X"E7", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FC", '1'),
      (X"9F23", X"F9", '1'),
      (X"9F23", X"F3", '1'),
      (X"9F23", X"E7", '1'),
      (X"9F23", X"CF", '1'),
      (X"9F23", X"9F", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"C3", '1'),
      (X"9F23", X"99", '1'),
      (X"9F23", X"91", '1'),
      (X"9F23", X"89", '1'),
      (X"9F23", X"99", '1'),
      (X"9F23", X"99", '1'),
      (X"9F23", X"C3", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"E7", '1'),
      (X"9F23", X"E7", '1'),
      (X"9F23", X"C7", '1'),
      (X"9F23", X"E7", '1'),
      (X"9F23", X"E7", '1'),
      (X"9F23", X"E7", '1'),
      (X"9F23", X"81", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"C3", '1'),
      (X"9F23", X"99", '1'),
      (X"9F23", X"F9", '1'),
      (X"9F23", X"F3", '1'),
      (X"9F23", X"CF", '1'),
      (X"9F23", X"9F", '1'),
      (X"9F23", X"81", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"C3", '1'),
      (X"9F23", X"99", '1'),
      (X"9F23", X"F9", '1'),
      (X"9F23", X"E3", '1'),
      (X"9F23", X"F9", '1'),
      (X"9F23", X"99", '1'),
      (X"9F23", X"C3", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"F9", '1'),
      (X"9F23", X"F1", '1'),
      (X"9F23", X"E1", '1'),
      (X"9F23", X"99", '1'),
      (X"9F23", X"80", '1'),
      (X"9F23", X"F9", '1'),
      (X"9F23", X"F9", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"81", '1'),
      (X"9F23", X"9F", '1'),
      (X"9F23", X"83", '1'),
      (X"9F23", X"F9", '1'),
      (X"9F23", X"F9", '1'),
      (X"9F23", X"99", '1'),
      (X"9F23", X"C3", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"C3", '1'),
      (X"9F23", X"99", '1'),
      (X"9F23", X"9F", '1'),
      (X"9F23", X"83", '1'),
      (X"9F23", X"99", '1'),
      (X"9F23", X"99", '1'),
      (X"9F23", X"C3", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"81", '1'),
      (X"9F23", X"99", '1'),
      (X"9F23", X"F3", '1'),
      (X"9F23", X"E7", '1'),
      (X"9F23", X"E7", '1'),
      (X"9F23", X"E7", '1'),
      (X"9F23", X"E7", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"C3", '1'),
      (X"9F23", X"99", '1'),
      (X"9F23", X"99", '1'),
      (X"9F23", X"C3", '1'),
      (X"9F23", X"99", '1'),
      (X"9F23", X"99", '1'),
      (X"9F23", X"C3", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"C3", '1'),
      (X"9F23", X"99", '1'),
      (X"9F23", X"99", '1'),
      (X"9F23", X"C1", '1'),
      (X"9F23", X"F9", '1'),
      (X"9F23", X"99", '1'),
      (X"9F23", X"C3", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"E7", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"E7", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"E7", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"E7", '1'),
      (X"9F23", X"E7", '1'),
      (X"9F23", X"CF", '1'),
      (X"9F23", X"F1", '1'),
      (X"9F23", X"E7", '1'),
      (X"9F23", X"CF", '1'),
      (X"9F23", X"9F", '1'),
      (X"9F23", X"CF", '1'),
      (X"9F23", X"E7", '1'),
      (X"9F23", X"F1", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"81", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"81", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"8F", '1'),
      (X"9F23", X"E7", '1'),
      (X"9F23", X"F3", '1'),
      (X"9F23", X"F9", '1'),
      (X"9F23", X"F3", '1'),
      (X"9F23", X"E7", '1'),
      (X"9F23", X"8F", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"C3", '1'),
      (X"9F23", X"99", '1'),
      (X"9F23", X"F9", '1'),
      (X"9F23", X"F3", '1'),
      (X"9F23", X"E7", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"E7", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'), -- 0x0FE00
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"F7", '1'),
      (X"9F23", X"E3", '1'),
      (X"9F23", X"C1", '1'),
      (X"9F23", X"80", '1'),
      (X"9F23", X"80", '1'),
      (X"9F23", X"E3", '1'),
      (X"9F23", X"C1", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"E7", '1'),
      (X"9F23", X"E7", '1'),
      (X"9F23", X"E7", '1'),
      (X"9F23", X"E7", '1'),
      (X"9F23", X"E7", '1'),
      (X"9F23", X"E7", '1'),
      (X"9F23", X"E7", '1'),
      (X"9F23", X"E7", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"CF", '1'),
      (X"9F23", X"CF", '1'),
      (X"9F23", X"CF", '1'),
      (X"9F23", X"CF", '1'),
      (X"9F23", X"CF", '1'),
      (X"9F23", X"CF", '1'),
      (X"9F23", X"CF", '1'),
      (X"9F23", X"CF", '1'),
      (X"9F23", X"F3", '1'),
      (X"9F23", X"F3", '1'),
      (X"9F23", X"F3", '1'),
      (X"9F23", X"F3", '1'),
      (X"9F23", X"F3", '1'),
      (X"9F23", X"F3", '1'),
      (X"9F23", X"F3", '1'),
      (X"9F23", X"F3", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"1F", '1'),
      (X"9F23", X"0F", '1'),
      (X"9F23", X"C7", '1'),
      (X"9F23", X"E7", '1'),
      (X"9F23", X"E7", '1'),
      (X"9F23", X"E7", '1'),
      (X"9F23", X"E7", '1'),
      (X"9F23", X"E3", '1'),
      (X"9F23", X"F0", '1'),
      (X"9F23", X"F8", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"E7", '1'),
      (X"9F23", X"E7", '1'),
      (X"9F23", X"C7", '1'),
      (X"9F23", X"0F", '1'),
      (X"9F23", X"1F", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"3F", '1'),
      (X"9F23", X"3F", '1'),
      (X"9F23", X"3F", '1'),
      (X"9F23", X"3F", '1'),
      (X"9F23", X"3F", '1'),
      (X"9F23", X"3F", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"3F", '1'),
      (X"9F23", X"1F", '1'),
      (X"9F23", X"8F", '1'),
      (X"9F23", X"C7", '1'),
      (X"9F23", X"E3", '1'),
      (X"9F23", X"F1", '1'),
      (X"9F23", X"F8", '1'),
      (X"9F23", X"FC", '1'),
      (X"9F23", X"FC", '1'),
      (X"9F23", X"F8", '1'),
      (X"9F23", X"F1", '1'),
      (X"9F23", X"E3", '1'),
      (X"9F23", X"C7", '1'),
      (X"9F23", X"8F", '1'),
      (X"9F23", X"1F", '1'),
      (X"9F23", X"3F", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"3F", '1'),
      (X"9F23", X"3F", '1'),
      (X"9F23", X"3F", '1'),
      (X"9F23", X"3F", '1'),
      (X"9F23", X"3F", '1'),
      (X"9F23", X"3F", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"FC", '1'),
      (X"9F23", X"FC", '1'),
      (X"9F23", X"FC", '1'),
      (X"9F23", X"FC", '1'),
      (X"9F23", X"FC", '1'),
      (X"9F23", X"FC", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"C3", '1'),
      (X"9F23", X"81", '1'),
      (X"9F23", X"81", '1'),
      (X"9F23", X"81", '1'),
      (X"9F23", X"81", '1'),
      (X"9F23", X"C3", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"C9", '1'),
      (X"9F23", X"80", '1'),
      (X"9F23", X"80", '1'),
      (X"9F23", X"80", '1'),
      (X"9F23", X"C1", '1'),
      (X"9F23", X"E3", '1'),
      (X"9F23", X"F7", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"9F", '1'),
      (X"9F23", X"9F", '1'),
      (X"9F23", X"9F", '1'),
      (X"9F23", X"9F", '1'),
      (X"9F23", X"9F", '1'),
      (X"9F23", X"9F", '1'),
      (X"9F23", X"9F", '1'),
      (X"9F23", X"9F", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"F8", '1'),
      (X"9F23", X"F0", '1'),
      (X"9F23", X"E3", '1'),
      (X"9F23", X"E7", '1'),
      (X"9F23", X"E7", '1'),
      (X"9F23", X"3C", '1'),
      (X"9F23", X"18", '1'),
      (X"9F23", X"81", '1'),
      (X"9F23", X"C3", '1'),
      (X"9F23", X"C3", '1'),
      (X"9F23", X"81", '1'),
      (X"9F23", X"18", '1'),
      (X"9F23", X"3C", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"C3", '1'),
      (X"9F23", X"81", '1'),
      (X"9F23", X"99", '1'),
      (X"9F23", X"99", '1'),
      (X"9F23", X"81", '1'),
      (X"9F23", X"C3", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"E7", '1'),
      (X"9F23", X"E7", '1'),
      (X"9F23", X"99", '1'),
      (X"9F23", X"99", '1'),
      (X"9F23", X"E7", '1'),
      (X"9F23", X"E7", '1'),
      (X"9F23", X"C3", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"F9", '1'),
      (X"9F23", X"F9", '1'),
      (X"9F23", X"F9", '1'),
      (X"9F23", X"F9", '1'),
      (X"9F23", X"F9", '1'),
      (X"9F23", X"F9", '1'),
      (X"9F23", X"F9", '1'),
      (X"9F23", X"F9", '1'),
      (X"9F23", X"F7", '1'),
      (X"9F23", X"E3", '1'),
      (X"9F23", X"C1", '1'),
      (X"9F23", X"80", '1'),
      (X"9F23", X"C1", '1'),
      (X"9F23", X"E3", '1'),
      (X"9F23", X"F7", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"E7", '1'),
      (X"9F23", X"E7", '1'),
      (X"9F23", X"E7", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"E7", '1'),
      (X"9F23", X"E7", '1'),
      (X"9F23", X"E7", '1'),
      (X"9F23", X"3F", '1'),
      (X"9F23", X"3F", '1'),
      (X"9F23", X"CF", '1'),
      (X"9F23", X"CF", '1'),
      (X"9F23", X"3F", '1'),
      (X"9F23", X"3F", '1'),
      (X"9F23", X"CF", '1'),
      (X"9F23", X"CF", '1'),
      (X"9F23", X"E7", '1'),
      (X"9F23", X"E7", '1'),
      (X"9F23", X"E7", '1'),
      (X"9F23", X"E7", '1'),
      (X"9F23", X"E7", '1'),
      (X"9F23", X"E7", '1'),
      (X"9F23", X"E7", '1'),
      (X"9F23", X"E7", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FC", '1'),
      (X"9F23", X"C1", '1'),
      (X"9F23", X"89", '1'),
      (X"9F23", X"C9", '1'),
      (X"9F23", X"C9", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"80", '1'),
      (X"9F23", X"C0", '1'),
      (X"9F23", X"E0", '1'),
      (X"9F23", X"F0", '1'),
      (X"9F23", X"F8", '1'),
      (X"9F23", X"FC", '1'),
      (X"9F23", X"FE", '1'),
      (X"9F23", X"FF", '1'), -- 0x0FF00
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"0F", '1'),
      (X"9F23", X"0F", '1'),
      (X"9F23", X"0F", '1'),
      (X"9F23", X"0F", '1'),
      (X"9F23", X"0F", '1'),
      (X"9F23", X"0F", '1'),
      (X"9F23", X"0F", '1'),
      (X"9F23", X"0F", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"3F", '1'),
      (X"9F23", X"3F", '1'),
      (X"9F23", X"3F", '1'),
      (X"9F23", X"3F", '1'),
      (X"9F23", X"3F", '1'),
      (X"9F23", X"3F", '1'),
      (X"9F23", X"3F", '1'),
      (X"9F23", X"3F", '1'),
      (X"9F23", X"33", '1'),
      (X"9F23", X"33", '1'),
      (X"9F23", X"CC", '1'),
      (X"9F23", X"CC", '1'),
      (X"9F23", X"33", '1'),
      (X"9F23", X"33", '1'),
      (X"9F23", X"CC", '1'),
      (X"9F23", X"CC", '1'),
      (X"9F23", X"FC", '1'),
      (X"9F23", X"FC", '1'),
      (X"9F23", X"FC", '1'),
      (X"9F23", X"FC", '1'),
      (X"9F23", X"FC", '1'),
      (X"9F23", X"FC", '1'),
      (X"9F23", X"FC", '1'),
      (X"9F23", X"FC", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"33", '1'),
      (X"9F23", X"33", '1'),
      (X"9F23", X"CC", '1'),
      (X"9F23", X"CC", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"01", '1'),
      (X"9F23", X"03", '1'),
      (X"9F23", X"07", '1'),
      (X"9F23", X"0F", '1'),
      (X"9F23", X"1F", '1'),
      (X"9F23", X"3F", '1'),
      (X"9F23", X"7F", '1'),
      (X"9F23", X"FC", '1'),
      (X"9F23", X"FC", '1'),
      (X"9F23", X"FC", '1'),
      (X"9F23", X"FC", '1'),
      (X"9F23", X"FC", '1'),
      (X"9F23", X"FC", '1'),
      (X"9F23", X"FC", '1'),
      (X"9F23", X"FC", '1'),
      (X"9F23", X"E7", '1'),
      (X"9F23", X"E7", '1'),
      (X"9F23", X"E7", '1'),
      (X"9F23", X"E0", '1'),
      (X"9F23", X"E0", '1'),
      (X"9F23", X"E7", '1'),
      (X"9F23", X"E7", '1'),
      (X"9F23", X"E7", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"F0", '1'),
      (X"9F23", X"F0", '1'),
      (X"9F23", X"F0", '1'),
      (X"9F23", X"F0", '1'),
      (X"9F23", X"E7", '1'),
      (X"9F23", X"E7", '1'),
      (X"9F23", X"E7", '1'),
      (X"9F23", X"E0", '1'),
      (X"9F23", X"E0", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"07", '1'),
      (X"9F23", X"07", '1'),
      (X"9F23", X"E7", '1'),
      (X"9F23", X"E7", '1'),
      (X"9F23", X"E7", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"E0", '1'),
      (X"9F23", X"E0", '1'),
      (X"9F23", X"E7", '1'),
      (X"9F23", X"E7", '1'),
      (X"9F23", X"E7", '1'),
      (X"9F23", X"E7", '1'),
      (X"9F23", X"E7", '1'),
      (X"9F23", X"E7", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"E7", '1'),
      (X"9F23", X"E7", '1'),
      (X"9F23", X"E7", '1'),
      (X"9F23", X"E7", '1'),
      (X"9F23", X"E7", '1'),
      (X"9F23", X"E7", '1'),
      (X"9F23", X"07", '1'),
      (X"9F23", X"07", '1'),
      (X"9F23", X"E7", '1'),
      (X"9F23", X"E7", '1'),
      (X"9F23", X"E7", '1'),
      (X"9F23", X"3F", '1'),
      (X"9F23", X"3F", '1'),
      (X"9F23", X"3F", '1'),
      (X"9F23", X"3F", '1'),
      (X"9F23", X"3F", '1'),
      (X"9F23", X"3F", '1'),
      (X"9F23", X"3F", '1'),
      (X"9F23", X"3F", '1'),
      (X"9F23", X"1F", '1'),
      (X"9F23", X"1F", '1'),
      (X"9F23", X"1F", '1'),
      (X"9F23", X"1F", '1'),
      (X"9F23", X"1F", '1'),
      (X"9F23", X"1F", '1'),
      (X"9F23", X"1F", '1'),
      (X"9F23", X"1F", '1'),
      (X"9F23", X"F8", '1'),
      (X"9F23", X"F8", '1'),
      (X"9F23", X"F8", '1'),
      (X"9F23", X"F8", '1'),
      (X"9F23", X"F8", '1'),
      (X"9F23", X"F8", '1'),
      (X"9F23", X"F8", '1'),
      (X"9F23", X"F8", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"FC", '1'),
      (X"9F23", X"FC", '1'),
      (X"9F23", X"FC", '1'),
      (X"9F23", X"FC", '1'),
      (X"9F23", X"FC", '1'),
      (X"9F23", X"FC", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"00", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"0F", '1'),
      (X"9F23", X"0F", '1'),
      (X"9F23", X"0F", '1'),
      (X"9F23", X"0F", '1'),
      (X"9F23", X"F0", '1'),
      (X"9F23", X"F0", '1'),
      (X"9F23", X"F0", '1'),
      (X"9F23", X"F0", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"E7", '1'),
      (X"9F23", X"E7", '1'),
      (X"9F23", X"E7", '1'),
      (X"9F23", X"07", '1'),
      (X"9F23", X"07", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"0F", '1'),
      (X"9F23", X"0F", '1'),
      (X"9F23", X"0F", '1'),
      (X"9F23", X"0F", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"FF", '1'),
      (X"9F23", X"0F", '1'),
      (X"9F23", X"0F", '1'),
      (X"9F23", X"0F", '1'),
      (X"9F23", X"0F", '1'),
      (X"9F23", X"F0", '1'),
      (X"9F23", X"F0", '1'),
      (X"9F23", X"F0", '1'),
      (X"9F23", X"F0", '1')
   );

   signal index : integer := 0;

begin

   -- This process generates the CPU accesses
   p_wr : process (clk_i)
   begin
      if rising_edge(clk_i) then
         wr_en_o <= '0';
         rd_en_o <= '0';
         if index < commands'length then
            addr_o    <= commands(index).addr(2 downto 0);
            if commands(index).wr_en = '1' then
               wr_en_o   <= '1';
               wr_data_o <= commands(index).data;
            else
               rd_en_o <= '1';
               exp_data_r <= commands(index).data;
            end if;
            index  <= index + 1;
         end if;
      end if;
   end process p_wr;

   -- This process verifies the result of the CPU reads.
   p_rd : process (clk_i)
   begin
      if rising_edge(clk_i) then
         if rd_en_o = '1' then
            assert rd_data_i = exp_data_r
               report "Read " & to_hstring(rd_data_i) & ", expected " & to_hstring(exp_data_r)
                  severity warning;
         end if;
      end if;
   end process p_rd;

end architecture structural;


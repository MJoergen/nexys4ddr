--------------------------------------
-- The Control Logic
--

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ctl is
   port (
      clk_i  : in  std_logic;
      rst_i  : in  std_logic;
      data_i : in  std_logic_vector( 7 downto 0);

      mem_rden_o      : out std_logic;                      -- Read from memory
      mem_wren_o      : out std_logic;                      -- Write to memory
      mem_addr_wren_o : out std_logic;                      -- Write to address hold register
      mem_addr_sel_o  : out std_logic_vector(3 downto 0);   -- Memory address select
      mem_data_sel_o  : out std_logic_vector(1 downto 0);   -- Memory data select
      reg_wren_o      : out std_logic;                      -- Write to register file
      reg_nr_o        : out std_logic_vector(1 downto 0);   -- Register number
      pc_sel_o        : out std_logic_vector(1 downto 0);   -- PC relect
      alu_func_o      : out std_logic_vector(3 downto 0);   -- ALU function
      clc_o           : out std_logic;                      -- Clear carry
      sr_alu_wren_o   : out std_logic;                      -- Write status register
      sp_sel_o        : out std_logic_vector(1 downto 0);   -- Stack pointer update

      debug_o : out std_logic_vector(10 downto 0)
   );
end ctl;

architecture Structural of ctl is

   signal cnt_r   : std_logic_vector(2 downto 0) := (others => '0');
   signal inst_r  : std_logic_vector(7 downto 0) := (others => '0');
   signal last    : std_logic;
   signal invalid : std_logic;

   signal ctl     : std_logic_vector(23 downto 0);

begin

   mem_rden_o      <= ctl(0);
   mem_wren_o      <= ctl(1);
   mem_addr_wren_o <= ctl(2);
   mem_addr_sel_o  <= ctl(6 downto 3);
   mem_data_sel_o  <= ctl(8 downto 7);
   reg_wren_o      <= ctl(9);
   reg_nr_o        <= ctl(11 downto 10);
   pc_sel_o        <= ctl(13 downto 12);
   sp_sel_o        <= ctl(15 downto 14);
   alu_func_o      <= ctl(19 downto 16);
   clc_o           <= ctl(20);
   sr_alu_wren_o   <= ctl(21);
   last            <= ctl(22);
   invalid         <= ctl(23);

   p_assert : process (clk_i)
   begin 
      if rising_edge(clk_i) then
         if rst_i = '0' then
            assert invalid = '0' report "Invalid opcode" severity failure;
         end if;
      end if;
   end process p_assert;

   debug_o( 7 downto 0) <= inst_r;
   debug_o(10 downto 8) <= cnt_r;

   -- Store the microinstruction counter
   p_cnt : process (clk_i)
   begin
      if rising_edge(clk_i) then
         cnt_r <= cnt_r + 1;

         if rst_i = '1' or last = '1' then
            cnt_r <= (others => '0');
         end if;
      end if;
   end process p_cnt;


   -- Store the current instruction
   p_inst : process (clk_i)
   begin
      if rising_edge(clk_i) then
         if cnt_r = 0 then
            inst_r <= data_i;
         end if;
      end if;
   end process p_inst;


   -- Combinatorial process
   process (cnt_r, inst_r)
   begin
      ctl <= B"0_0_0_0_0000_00_00_00_0_00_0000_0_0_0";  -- Default value to avoid latch.

      if cnt_r = 0 then
         ctl <= B"0_0_0_0_0000_00_00_00_0_00_0000_0_0_1";  -- Default value to avoid latch.
      end if;

      if cnt_r = 1 then
         case inst_r is
            when X"00" => ctl <= B"0_0_0_0_0000_10_11_00_0_01_0010_0_1_0"; -- BRK b
            when X"01" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ORA (d,X)
            when X"02" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"03" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"04" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"05" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ORA d
            when X"06" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ASL d
            when X"07" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"08" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- PHP
            when X"09" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ORA #
            when X"0A" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ASL A
            when X"0B" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"0C" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"0D" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ORA a
            when X"0E" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ASL a
            when X"0F" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";

            when X"10" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- BPL r
            when X"11" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ORA (d),Y
            when X"12" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"13" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"14" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"15" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ORA d,X
            when X"16" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ASL d,X
            when X"17" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"18" => ctl <= B"0_1_0_1_0000_00_11_00_0_00_0000_0_0_0"; -- CLC
            when X"19" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ORA a,Y
            when X"1A" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"1B" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"1C" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"1D" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ORA a,X
            when X"1E" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ASL a,X
            when X"1F" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";

            when X"20" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- JSR a
            when X"21" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- AND (d,X)
            when X"22" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"23" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"24" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- BIT d
            when X"25" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- AND d
            when X"26" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ROL d
            when X"27" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"28" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- PLP
            when X"29" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- AND #
            when X"2A" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ROL A
            when X"2B" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"2C" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- BIT a
            when X"2D" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- AND a
            when X"2E" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ROL a
            when X"2F" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";

            when X"30" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- BMI r
            when X"31" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- AND (d),Y
            when X"32" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"33" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"34" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"35" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- AND d,X
            when X"36" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ROL d,X
            when X"37" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"38" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- SEC
            when X"39" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- AND a,Y
            when X"3A" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"3B" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"3C" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"3D" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- AND a,X
            when X"3E" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ROL a,X
            when X"3F" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";

            when X"40" => ctl <= B"0_0_0_0_0000_01_11_00_0_00_0000_0_0_0"; -- RTI
            when X"41" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- EOR (d,X)
            when X"42" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"43" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"44" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"45" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- EOR d
            when X"46" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LSR d
            when X"47" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"48" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- PHA
            when X"49" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- EOR #
            when X"4A" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LSR A
            when X"4B" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"4C" => ctl <= B"0_0_0_0_0000_00_00_00_0_00_0000_1_0_1"; -- JMP a
            when X"4D" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- EOR a
            when X"4E" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LSR a
            when X"4F" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";

            when X"50" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- BVC r
            when X"51" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- EOR (d),Y
            when X"52" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"53" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"54" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"55" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- EOR d,X
            when X"56" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LSR d,X
            when X"57" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"58" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- CLI
            when X"59" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- EOR a,Y
            when X"5A" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"5B" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"5C" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"5D" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- EOR a,X
            when X"5E" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LSR a,X
            when X"5F" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";

            when X"60" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- RTS
            when X"61" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ADC (d,X)
            when X"62" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"63" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"64" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"65" => ctl <= B"0_0_0_0_0000_00_00_00_0_00_0000_1_0_1"; -- ADC d
            when X"66" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ROR d
            when X"67" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"68" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- PLA
            when X"69" => ctl <= B"0_1_1_0_0011_00_00_00_1_00_0000_0_0_1"; -- ADC #
            when X"6A" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ROR A
            when X"6B" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"6C" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- JMP (a)
            when X"6D" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ADC a
            when X"6E" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ROR a
            when X"6F" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";

            when X"70" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- BVS r
            when X"71" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ADC (d),Y
            when X"72" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"73" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"74" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"75" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ADC d,X
            when X"76" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ROR d,X
            when X"77" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"78" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- SEI
            when X"79" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ADC a,Y
            when X"7A" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"7B" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"7C" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"7D" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ADC a,X
            when X"7E" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ROR a,X
            when X"7F" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";

            when X"80" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"81" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- STA (d,X)
            when X"82" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"83" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"84" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- STY
            when X"85" => ctl <= B"0_0_0_0_0000_00_00_00_0_00_0000_1_0_1"; -- STA d
            when X"86" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- STX d
            when X"87" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"88" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- DEY
            when X"89" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"8A" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- TXA
            when X"8B" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; 
            when X"8C" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- STY a
            when X"8D" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- STA a
            when X"8E" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- STX a
            when X"8F" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";

            when X"90" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- BCC r
            when X"91" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- STA (d),Y
            when X"92" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"93" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"94" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- STY d,X
            when X"95" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- STA d,X
            when X"96" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- STX d,Y
            when X"97" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"98" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- TYA
            when X"99" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- STA a,Y
            when X"9A" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- TXS
            when X"9B" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"9C" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"9D" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- STA a,X
            when X"9E" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"9F" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";

            when X"A0" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LDY #
            when X"A1" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LDA (d,X)
            when X"A2" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LDX #
            when X"A3" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"A4" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LDY d
            when X"A5" => ctl <= B"0_0_0_0_0000_00_00_00_0_00_0000_1_0_1"; -- LDA d
            when X"A6" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LDX d
            when X"A7" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"A8" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- TAY
            when X"A9" => ctl <= B"0_1_0_0_0101_00_00_00_1_00_0000_0_0_1"; -- LDA #
            when X"AA" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- TAX
            when X"AB" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"AC" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LDY a
            when X"AD" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LDA a
            when X"AE" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LDX a
            when X"AF" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";

            when X"B0" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- BCS r
            when X"B1" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LDA (d),Y
            when X"B2" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"B3" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"B4" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LDY d,X
            when X"B5" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LDA d,X
            when X"B6" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LDX d,Y
            when X"B7" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"B8" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- CLV
            when X"B9" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LDA a,Y
            when X"BA" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- TSX
            when X"BB" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"BC" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LDY a,X
            when X"BD" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LDA a,X
            when X"BE" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LDX a,Y
            when X"BF" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";

            when X"C0" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- CPY #
            when X"C1" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- CMP (d,X)
            when X"C2" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"C3" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"C4" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- CPY d
            when X"C5" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- CMP d
            when X"C6" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- DEC d
            when X"C7" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"C8" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- INY
            when X"C9" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- CMP #
            when X"CA" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- DEX
            when X"CB" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"CC" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- CPY a
            when X"CD" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- CMP a
            when X"CE" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- DEC a
            when X"CF" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";

            when X"D0" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- BNE r
            when X"D1" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- CMP (d),Y
            when X"D2" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"D3" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"D4" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"D5" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- CMP d,X
            when X"D6" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- DEC d,X
            when X"D7" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"D8" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- CLD
            when X"D9" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- CMP a,Y
            when X"DA" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"DB" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"DC" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"DD" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- CMP a,X
            when X"DE" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- DEC a,X
            when X"DF" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";

            when X"E0" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- CPX #
            when X"E1" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- SBC (d,X)
            when X"E2" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"E3" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"E4" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- CPX d
            when X"E5" => ctl <= B"0_0_0_0_0000_00_00_00_0_00_0000_1_0_1"; -- SBC d
            when X"E6" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- INC d
            when X"E7" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"E8" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- INX
            when X"E9" => ctl <= B"0_1_1_0_0111_00_00_00_1_00_0000_0_0_1"; -- SBC #
            when X"EA" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- NOP
            when X"EB" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"EC" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- CPX a
            when X"ED" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- SBC a
            when X"EE" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- INC a
            when X"EF" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";

            when X"F0" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- BEQ r
            when X"F1" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- SBC (d),Y
            when X"F2" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"F3" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"F4" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"F5" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- SBC d,X
            when X"F6" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- INC d,X
            when X"F7" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"F8" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- SED
            when X"F9" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- SBC a,Y
            when X"FA" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"FB" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"FC" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"FD" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- SBC a,X
            when X"FE" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- INC a,X
            when X"FF" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";

            when others =>ctl <= B"0_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; 
         end case;
      end if;

      if cnt_r = 2 then
         case inst_r is
            when X"00" => ctl <= B"0_0_0_0_0000_10_11_00_0_10_0010_0_1_0"; -- BRK b
            when X"01" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ORA (d,X)
            when X"02" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"03" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"04" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"05" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ORA d
            when X"06" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ASL d
            when X"07" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"08" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- PHP
            when X"09" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ORA #
            when X"0A" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ASL A
            when X"0B" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"0C" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"0D" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ORA a
            when X"0E" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ASL a
            when X"0F" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";

            when X"10" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- BPL r
            when X"11" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ORA (d),Y
            when X"12" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"13" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"14" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"15" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ORA d,X
            when X"16" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ASL d,X
            when X"17" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"18" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- CLC
            when X"19" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ORA a,Y
            when X"1A" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"1B" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"1C" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"1D" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ORA a,X
            when X"1E" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ASL a,X
            when X"1F" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";

            when X"20" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- JSR a
            when X"21" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- AND (d,X)
            when X"22" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"23" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"24" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- BIT d
            when X"25" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- AND d
            when X"26" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ROL d
            when X"27" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"28" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- PLP
            when X"29" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- AND #
            when X"2A" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ROL A
            when X"2B" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"2C" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- BIT a
            when X"2D" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- AND a
            when X"2E" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ROL a
            when X"2F" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";

            when X"30" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- BMI r
            when X"31" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- AND (d),Y
            when X"32" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"33" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"34" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"35" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- AND d,X
            when X"36" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ROL d,X
            when X"37" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"38" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- SEC
            when X"39" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- AND a,Y
            when X"3A" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"3B" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"3C" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"3D" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- AND a,X
            when X"3E" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ROL a,X
            when X"3F" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";

            when X"40" => ctl <= B"0_0_0_0_0000_01_11_00_0_00_0010_0_0_1"; -- RTI
            when X"41" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- EOR (d,X)
            when X"42" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"43" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"44" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"45" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- EOR d
            when X"46" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LSR d
            when X"47" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"48" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- PHA
            when X"49" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- EOR #
            when X"4A" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LSR A
            when X"4B" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"4C" => ctl <= B"0_1_0_0_0000_00_01_00_0_00_0000_0_0_1"; -- JMP a
            when X"4D" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- EOR a
            when X"4E" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LSR a
            when X"4F" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";

            when X"50" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- BVC r
            when X"51" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- EOR (d),Y
            when X"52" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"53" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"54" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"55" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- EOR d,X
            when X"56" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LSR d,X
            when X"57" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"58" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- CLI
            when X"59" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- EOR a,Y
            when X"5A" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"5B" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"5C" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"5D" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- EOR a,X
            when X"5E" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LSR a,X
            when X"5F" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";

            when X"60" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- RTS
            when X"61" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ADC (d,X)
            when X"62" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"63" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"64" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"65" => ctl <= B"0_1_1_0_0011_00_11_00_1_00_0001_0_0_1"; -- ADC d
            when X"66" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ROR d
            when X"67" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"68" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- PLA
            when X"69" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ADC #
            when X"6A" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ROR A
            when X"6B" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"6C" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- JMP (a)
            when X"6D" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ADC a
            when X"6E" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ROR a
            when X"6F" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";

            when X"70" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- BVS r
            when X"71" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ADC (d),Y
            when X"72" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"73" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"74" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"75" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ADC d,X
            when X"76" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ROR d,X
            when X"77" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"78" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- SEI
            when X"79" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ADC a,Y
            when X"7A" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"7B" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"7C" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"7D" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ADC a,X
            when X"7E" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ROR a,X
            when X"7F" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";

            when X"80" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"81" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- STA (d,X)
            when X"82" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"83" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"84" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- STY
            when X"85" => ctl <= B"0_1_0_0_0000_00_11_00_0_00_0001_0_1_0"; -- STA d
            when X"86" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- STX d
            when X"87" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"88" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- DEY
            when X"89" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"8A" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- TXA
            when X"8B" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; 
            when X"8C" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- STY a
            when X"8D" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- STA a
            when X"8E" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- STX a
            when X"8F" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";

            when X"90" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- BCC r
            when X"91" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- STA (d),Y
            when X"92" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"93" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"94" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- STY d,X
            when X"95" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- STA d,X
            when X"96" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- STX d,Y
            when X"97" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"98" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- TYA
            when X"99" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- STA a,Y
            when X"9A" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- TXS
            when X"9B" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"9C" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"9D" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- STA a,X
            when X"9E" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"9F" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";

            when X"A0" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LDY #
            when X"A1" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LDA (d,X)
            when X"A2" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LDX #
            when X"A3" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"A4" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LDY d
            when X"A5" => ctl <= B"0_1_0_0_0101_00_11_00_1_00_0001_0_0_1"; -- LDA d
            when X"A6" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LDX d
            when X"A7" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"A8" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- TAY
            when X"A9" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LDA #
            when X"AA" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- TAX
            when X"AB" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"AC" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LDY a
            when X"AD" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LDA a
            when X"AE" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LDX a
            when X"AF" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";

            when X"B0" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- BCS r
            when X"B1" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LDA (d),Y
            when X"B2" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"B3" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"B4" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LDY d,X
            when X"B5" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LDA d,X
            when X"B6" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LDX d,Y
            when X"B7" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"B8" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- CLV
            when X"B9" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LDA a,Y
            when X"BA" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- TSX
            when X"BB" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"BC" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LDY a,X
            when X"BD" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LDA a,X
            when X"BE" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LDX a,Y
            when X"BF" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";

            when X"C0" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- CPY #
            when X"C1" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- CMP (d,X)
            when X"C2" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"C3" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"C4" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- CPY d
            when X"C5" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- CMP d
            when X"C6" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- DEC d
            when X"C7" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"C8" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- INY
            when X"C9" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- CMP #
            when X"CA" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- DEX
            when X"CB" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"CC" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- CPY a
            when X"CD" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- CMP a
            when X"CE" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- DEC a
            when X"CF" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";

            when X"D0" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- BNE r
            when X"D1" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- CMP (d),Y
            when X"D2" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"D3" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"D4" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"D5" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- CMP d,X
            when X"D6" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- DEC d,X
            when X"D7" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"D8" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- CLD
            when X"D9" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- CMP a,Y
            when X"DA" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"DB" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"DC" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"DD" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- CMP a,X
            when X"DE" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- DEC a,X
            when X"DF" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";

            when X"E0" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- CPX #
            when X"E1" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- SBC (d,X)
            when X"E2" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"E3" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"E4" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- CPX d
            when X"E5" => ctl <= B"0_1_1_0_0111_00_11_00_1_00_0001_0_0_1"; -- SBC d
            when X"E6" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- INC d
            when X"E7" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"E8" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- INX
            when X"E9" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- SBC #
            when X"EA" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- NOP
            when X"EB" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"EC" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- CPX a
            when X"ED" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- SBC a
            when X"EE" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- INC a
            when X"EF" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";

            when X"F0" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- BEQ r
            when X"F1" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- SBC (d),Y
            when X"F2" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"F3" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"F4" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"F5" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- SBC d,X
            when X"F6" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- INC d,X
            when X"F7" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"F8" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- SED
            when X"F9" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- SBC a,Y
            when X"FA" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"FB" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"FC" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"FD" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- SBC a,X
            when X"FE" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- INC a,X
            when X"FF" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";

            when others =>ctl <= B"0_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; 
         end case;
      end if;

      if cnt_r = 3 then
         case inst_r is
            when X"00" => ctl <= B"0_0_0_0_0000_10_11_00_0_11_0010_0_1_0"; -- BRK b
            when X"01" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ORA (d,X)
            when X"02" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"03" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"04" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"05" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ORA d
            when X"06" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ASL d
            when X"07" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"08" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- PHP
            when X"09" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ORA #
            when X"0A" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ASL A
            when X"0B" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"0C" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"0D" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ORA a
            when X"0E" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ASL a
            when X"0F" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";

            when X"10" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- BPL r
            when X"11" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ORA (d),Y
            when X"12" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"13" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"14" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"15" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ORA d,X
            when X"16" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ASL d,X
            when X"17" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"18" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- CLC
            when X"19" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ORA a,Y
            when X"1A" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"1B" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"1C" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"1D" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ORA a,X
            when X"1E" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ASL a,X
            when X"1F" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";

            when X"20" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- JSR a
            when X"21" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- AND (d,X)
            when X"22" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"23" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"24" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- BIT d
            when X"25" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- AND d
            when X"26" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ROL d
            when X"27" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"28" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- PLP
            when X"29" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- AND #
            when X"2A" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ROL A
            when X"2B" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"2C" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- BIT a
            when X"2D" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- AND a
            when X"2E" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ROL a
            when X"2F" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";

            when X"30" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- BMI r
            when X"31" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- AND (d),Y
            when X"32" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"33" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"34" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"35" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- AND d,X
            when X"36" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ROL d,X
            when X"37" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"38" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- SEC
            when X"39" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- AND a,Y
            when X"3A" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"3B" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"3C" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"3D" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- AND a,X
            when X"3E" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ROL a,X
            when X"3F" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";

            when X"40" => ctl <= B"0_0_0_0_0000_01_11_00_0_00_0010_1_0_1"; -- RTI
            when X"41" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- EOR (d,X)
            when X"42" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"43" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"44" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"45" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- EOR d
            when X"46" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LSR d
            when X"47" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"48" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- PHA
            when X"49" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- EOR #
            when X"4A" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LSR A
            when X"4B" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"4C" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- JMP a
            when X"4D" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- EOR a
            when X"4E" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LSR a
            when X"4F" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";

            when X"50" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- BVC r
            when X"51" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- EOR (d),Y
            when X"52" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"53" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"54" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"55" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- EOR d,X
            when X"56" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LSR d,X
            when X"57" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"58" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- CLI
            when X"59" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- EOR a,Y
            when X"5A" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"5B" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"5C" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"5D" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- EOR a,X
            when X"5E" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LSR a,X
            when X"5F" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";

            when X"60" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- RTS
            when X"61" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ADC (d,X)
            when X"62" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"63" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"64" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"65" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ADC d
            when X"66" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ROR d
            when X"67" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"68" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- PLA
            when X"69" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ADC #
            when X"6A" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ROR A
            when X"6B" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"6C" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- JMP (a)
            when X"6D" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ADC a
            when X"6E" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ROR a
            when X"6F" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";

            when X"70" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- BVS r
            when X"71" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ADC (d),Y
            when X"72" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"73" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"74" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"75" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ADC d,X
            when X"76" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ROR d,X
            when X"77" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"78" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- SEI
            when X"79" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ADC a,Y
            when X"7A" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"7B" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"7C" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"7D" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ADC a,X
            when X"7E" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ROR a,X
            when X"7F" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";

            when X"80" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"81" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- STA (d,X)
            when X"82" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"83" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"84" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- STY
            when X"85" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- STA d
            when X"86" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- STX d
            when X"87" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"88" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- DEY
            when X"89" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"8A" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- TXA
            when X"8B" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; 
            when X"8C" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- STY a
            when X"8D" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- STA a
            when X"8E" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- STX a
            when X"8F" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";

            when X"90" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- BCC r
            when X"91" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- STA (d),Y
            when X"92" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"93" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"94" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- STY d,X
            when X"95" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- STA d,X
            when X"96" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- STX d,Y
            when X"97" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"98" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- TYA
            when X"99" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- STA a,Y
            when X"9A" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- TXS
            when X"9B" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"9C" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"9D" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- STA a,X
            when X"9E" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"9F" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";

            when X"A0" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LDY #
            when X"A1" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LDA (d,X)
            when X"A2" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LDX #
            when X"A3" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"A4" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LDY d
            when X"A5" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LDA d
            when X"A6" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LDX d
            when X"A7" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"A8" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- TAY
            when X"A9" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LDA #
            when X"AA" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- TAX
            when X"AB" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"AC" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LDY a
            when X"AD" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LDA a
            when X"AE" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LDX a
            when X"AF" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";

            when X"B0" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- BCS r
            when X"B1" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LDA (d),Y
            when X"B2" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"B3" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"B4" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LDY d,X
            when X"B5" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LDA d,X
            when X"B6" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LDX d,Y
            when X"B7" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"B8" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- CLV
            when X"B9" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LDA a,Y
            when X"BA" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- TSX
            when X"BB" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"BC" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LDY a,X
            when X"BD" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LDA a,X
            when X"BE" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LDX a,Y
            when X"BF" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";

            when X"C0" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- CPY #
            when X"C1" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- CMP (d,X)
            when X"C2" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"C3" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"C4" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- CPY d
            when X"C5" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- CMP d
            when X"C6" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- DEC d
            when X"C7" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"C8" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- INY
            when X"C9" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- CMP #
            when X"CA" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- DEX
            when X"CB" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"CC" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- CPY a
            when X"CD" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- CMP a
            when X"CE" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- DEC a
            when X"CF" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";

            when X"D0" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- BNE r
            when X"D1" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- CMP (d),Y
            when X"D2" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"D3" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"D4" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"D5" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- CMP d,X
            when X"D6" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- DEC d,X
            when X"D7" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"D8" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- CLD
            when X"D9" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- CMP a,Y
            when X"DA" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"DB" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"DC" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"DD" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- CMP a,X
            when X"DE" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- DEC a,X
            when X"DF" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";

            when X"E0" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- CPX #
            when X"E1" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- SBC (d,X)
            when X"E2" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"E3" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"E4" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- CPX d
            when X"E5" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- SBC d
            when X"E6" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- INC d
            when X"E7" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"E8" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- INX
            when X"E9" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- SBC #
            when X"EA" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- NOP
            when X"EB" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"EC" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- CPX a
            when X"ED" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- SBC a
            when X"EE" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- INC a
            when X"EF" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";

            when X"F0" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- BEQ r
            when X"F1" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- SBC (d),Y
            when X"F2" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"F3" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"F4" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"F5" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- SBC d,X
            when X"F6" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- INC d,X
            when X"F7" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"F8" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- SED
            when X"F9" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- SBC a,Y
            when X"FA" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"FB" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"FC" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"FD" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- SBC a,X
            when X"FE" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- INC a,X
            when X"FF" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";

            when others =>ctl <= B"0_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; 
         end case;
      end if;

      if cnt_r = 4 then
         case inst_r is
            when X"00" => ctl <= B"0_0_0_0_0000_00_11_00_0_00_1110_1_0_1"; -- BRK b
            when X"01" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ORA (d,X)
            when X"02" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"03" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"04" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"05" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ORA d
            when X"06" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ASL d
            when X"07" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"08" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- PHP
            when X"09" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ORA #
            when X"0A" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ASL A
            when X"0B" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"0C" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"0D" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ORA a
            when X"0E" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ASL a
            when X"0F" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";

            when X"10" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- BPL r
            when X"11" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ORA (d),Y
            when X"12" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"13" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"14" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"15" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ORA d,X
            when X"16" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ASL d,X
            when X"17" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"18" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- CLC
            when X"19" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ORA a,Y
            when X"1A" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"1B" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"1C" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"1D" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ORA a,X
            when X"1E" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ASL a,X
            when X"1F" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";

            when X"20" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- JSR a
            when X"21" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- AND (d,X)
            when X"22" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"23" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"24" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- BIT d
            when X"25" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- AND d
            when X"26" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ROL d
            when X"27" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"28" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- PLP
            when X"29" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- AND #
            when X"2A" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ROL A
            when X"2B" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"2C" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- BIT a
            when X"2D" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- AND a
            when X"2E" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ROL a
            when X"2F" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";

            when X"30" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- BMI r
            when X"31" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- AND (d),Y
            when X"32" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"33" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"34" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"35" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- AND d,X
            when X"36" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ROL d,X
            when X"37" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"38" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- SEC
            when X"39" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- AND a,Y
            when X"3A" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"3B" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"3C" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"3D" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- AND a,X
            when X"3E" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ROL a,X
            when X"3F" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";

            when X"40" => ctl <= B"0_1_0_0_0000_00_01_00_0_00_0000_0_0_0"; -- RTI
            when X"41" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- EOR (d,X)
            when X"42" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"43" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"44" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"45" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- EOR d
            when X"46" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LSR d
            when X"47" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"48" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- PHA
            when X"49" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- EOR #
            when X"4A" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LSR A
            when X"4B" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"4C" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- JMP a
            when X"4D" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- EOR a
            when X"4E" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LSR a
            when X"4F" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";

            when X"50" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- BVC r
            when X"51" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- EOR (d),Y
            when X"52" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"53" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"54" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"55" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- EOR d,X
            when X"56" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LSR d,X
            when X"57" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"58" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- CLI
            when X"59" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- EOR a,Y
            when X"5A" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"5B" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"5C" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"5D" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- EOR a,X
            when X"5E" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LSR a,X
            when X"5F" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";

            when X"60" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- RTS
            when X"61" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ADC (d,X)
            when X"62" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"63" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"64" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"65" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ADC d
            when X"66" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ROR d
            when X"67" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"68" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- PLA
            when X"69" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ADC #
            when X"6A" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ROR A
            when X"6B" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"6C" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- JMP (a)
            when X"6D" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ADC a
            when X"6E" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ROR a
            when X"6F" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";

            when X"70" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- BVS r
            when X"71" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ADC (d),Y
            when X"72" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"73" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"74" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"75" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ADC d,X
            when X"76" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ROR d,X
            when X"77" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"78" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- SEI
            when X"79" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ADC a,Y
            when X"7A" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"7B" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"7C" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"7D" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ADC a,X
            when X"7E" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ROR a,X
            when X"7F" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";

            when X"80" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"81" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- STA (d,X)
            when X"82" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"83" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"84" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- STY
            when X"85" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- STA d
            when X"86" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- STX d
            when X"87" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"88" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- DEY
            when X"89" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"8A" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- TXA
            when X"8B" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; 
            when X"8C" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- STY a
            when X"8D" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- STA a
            when X"8E" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- STX a
            when X"8F" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";

            when X"90" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- BCC r
            when X"91" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- STA (d),Y
            when X"92" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"93" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"94" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- STY d,X
            when X"95" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- STA d,X
            when X"96" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- STX d,Y
            when X"97" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"98" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- TYA
            when X"99" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- STA a,Y
            when X"9A" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- TXS
            when X"9B" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"9C" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"9D" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- STA a,X
            when X"9E" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"9F" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";

            when X"A0" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LDY #
            when X"A1" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LDA (d,X)
            when X"A2" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LDX #
            when X"A3" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"A4" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LDY d
            when X"A5" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LDA d
            when X"A6" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LDX d
            when X"A7" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"A8" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- TAY
            when X"A9" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LDA #
            when X"AA" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- TAX
            when X"AB" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"AC" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LDY a
            when X"AD" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LDA a
            when X"AE" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LDX a
            when X"AF" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";

            when X"B0" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- BCS r
            when X"B1" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LDA (d),Y
            when X"B2" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"B3" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"B4" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LDY d,X
            when X"B5" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LDA d,X
            when X"B6" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LDX d,Y
            when X"B7" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"B8" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- CLV
            when X"B9" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LDA a,Y
            when X"BA" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- TSX
            when X"BB" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"BC" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LDY a,X
            when X"BD" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LDA a,X
            when X"BE" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LDX a,Y
            when X"BF" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";

            when X"C0" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- CPY #
            when X"C1" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- CMP (d,X)
            when X"C2" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"C3" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"C4" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- CPY d
            when X"C5" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- CMP d
            when X"C6" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- DEC d
            when X"C7" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"C8" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- INY
            when X"C9" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- CMP #
            when X"CA" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- DEX
            when X"CB" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"CC" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- CPY a
            when X"CD" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- CMP a
            when X"CE" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- DEC a
            when X"CF" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";

            when X"D0" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- BNE r
            when X"D1" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- CMP (d),Y
            when X"D2" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"D3" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"D4" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"D5" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- CMP d,X
            when X"D6" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- DEC d,X
            when X"D7" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"D8" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- CLD
            when X"D9" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- CMP a,Y
            when X"DA" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"DB" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"DC" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"DD" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- CMP a,X
            when X"DE" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- DEC a,X
            when X"DF" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";

            when X"E0" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- CPX #
            when X"E1" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- SBC (d,X)
            when X"E2" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"E3" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"E4" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- CPX d
            when X"E5" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- SBC d
            when X"E6" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- INC d
            when X"E7" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"E8" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- INX
            when X"E9" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- SBC #
            when X"EA" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- NOP
            when X"EB" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"EC" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- CPX a
            when X"ED" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- SBC a
            when X"EE" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- INC a
            when X"EF" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";

            when X"F0" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- BEQ r
            when X"F1" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- SBC (d),Y
            when X"F2" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"F3" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"F4" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"F5" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- SBC d,X
            when X"F6" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- INC d,X
            when X"F7" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"F8" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- SED
            when X"F9" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- SBC a,Y
            when X"FA" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"FB" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"FC" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"FD" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- SBC a,X
            when X"FE" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- INC a,X
            when X"FF" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";

            when others =>ctl <= B"0_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; 
         end case;
      end if;

      if cnt_r = 5 then
         case inst_r is
            when X"00" => ctl <= B"0_1_0_0_0000_00_01_00_0_00_1111_0_0_1"; -- BRK b
            when X"01" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ORA (d,X)
            when X"02" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"03" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"04" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"05" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ORA d
            when X"06" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ASL d
            when X"07" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"08" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- PHP
            when X"09" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ORA #
            when X"0A" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ASL A
            when X"0B" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"0C" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"0D" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ORA a
            when X"0E" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ASL a
            when X"0F" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";

            when X"10" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- BPL r
            when X"11" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ORA (d),Y
            when X"12" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"13" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"14" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"15" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ORA d,X
            when X"16" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ASL d,X
            when X"17" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"18" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- CLC
            when X"19" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ORA a,Y
            when X"1A" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"1B" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"1C" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"1D" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ORA a,X
            when X"1E" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ASL a,X
            when X"1F" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";

            when X"20" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- JSR a
            when X"21" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- AND (d,X)
            when X"22" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"23" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"24" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- BIT d
            when X"25" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- AND d
            when X"26" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ROL d
            when X"27" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"28" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- PLP
            when X"29" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- AND #
            when X"2A" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ROL A
            when X"2B" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"2C" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- BIT a
            when X"2D" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- AND a
            when X"2E" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ROL a
            when X"2F" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";

            when X"30" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- BMI r
            when X"31" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- AND (d),Y
            when X"32" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"33" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"34" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"35" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- AND d,X
            when X"36" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ROL d,X
            when X"37" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"38" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- SEC
            when X"39" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- AND a,Y
            when X"3A" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"3B" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"3C" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"3D" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- AND a,X
            when X"3E" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ROL a,X
            when X"3F" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";

            when X"40" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- RTI
            when X"41" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- EOR (d,X)
            when X"42" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"43" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"44" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"45" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- EOR d
            when X"46" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LSR d
            when X"47" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"48" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- PHA
            when X"49" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- EOR #
            when X"4A" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LSR A
            when X"4B" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"4C" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- JMP a
            when X"4D" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- EOR a
            when X"4E" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LSR a
            when X"4F" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";

            when X"50" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- BVC r
            when X"51" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- EOR (d),Y
            when X"52" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"53" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"54" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"55" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- EOR d,X
            when X"56" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LSR d,X
            when X"57" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"58" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- CLI
            when X"59" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- EOR a,Y
            when X"5A" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"5B" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"5C" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"5D" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- EOR a,X
            when X"5E" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LSR a,X
            when X"5F" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";

            when X"60" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- RTS
            when X"61" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ADC (d,X)
            when X"62" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"63" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"64" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"65" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ADC d
            when X"66" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ROR d
            when X"67" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"68" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- PLA
            when X"69" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ADC #
            when X"6A" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ROR A
            when X"6B" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"6C" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- JMP (a)
            when X"6D" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ADC a
            when X"6E" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ROR a
            when X"6F" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";

            when X"70" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- BVS r
            when X"71" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ADC (d),Y
            when X"72" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"73" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"74" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"75" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ADC d,X
            when X"76" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ROR d,X
            when X"77" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"78" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- SEI
            when X"79" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ADC a,Y
            when X"7A" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"7B" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"7C" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"7D" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ADC a,X
            when X"7E" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ROR a,X
            when X"7F" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";

            when X"80" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"81" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- STA (d,X)
            when X"82" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"83" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"84" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- STY
            when X"85" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- STA d
            when X"86" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- STX d
            when X"87" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"88" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- DEY
            when X"89" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"8A" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- TXA
            when X"8B" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; 
            when X"8C" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- STY a
            when X"8D" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- STA a
            when X"8E" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- STX a
            when X"8F" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";

            when X"90" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- BCC r
            when X"91" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- STA (d),Y
            when X"92" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"93" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"94" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- STY d,X
            when X"95" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- STA d,X
            when X"96" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- STX d,Y
            when X"97" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"98" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- TYA
            when X"99" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- STA a,Y
            when X"9A" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- TXS
            when X"9B" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"9C" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"9D" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- STA a,X
            when X"9E" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"9F" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";

            when X"A0" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LDY #
            when X"A1" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LDA (d,X)
            when X"A2" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LDX #
            when X"A3" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"A4" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LDY d
            when X"A5" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LDA d
            when X"A6" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LDX d
            when X"A7" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"A8" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- TAY
            when X"A9" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LDA #
            when X"AA" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- TAX
            when X"AB" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"AC" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LDY a
            when X"AD" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LDA a
            when X"AE" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LDX a
            when X"AF" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";

            when X"B0" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- BCS r
            when X"B1" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LDA (d),Y
            when X"B2" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"B3" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"B4" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LDY d,X
            when X"B5" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LDA d,X
            when X"B6" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LDX d,Y
            when X"B7" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"B8" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- CLV
            when X"B9" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LDA a,Y
            when X"BA" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- TSX
            when X"BB" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"BC" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LDY a,X
            when X"BD" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LDA a,X
            when X"BE" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LDX a,Y
            when X"BF" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";

            when X"C0" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- CPY #
            when X"C1" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- CMP (d,X)
            when X"C2" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"C3" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"C4" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- CPY d
            when X"C5" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- CMP d
            when X"C6" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- DEC d
            when X"C7" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"C8" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- INY
            when X"C9" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- CMP #
            when X"CA" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- DEX
            when X"CB" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"CC" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- CPY a
            when X"CD" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- CMP a
            when X"CE" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- DEC a
            when X"CF" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";

            when X"D0" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- BNE r
            when X"D1" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- CMP (d),Y
            when X"D2" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"D3" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"D4" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"D5" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- CMP d,X
            when X"D6" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- DEC d,X
            when X"D7" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"D8" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- CLD
            when X"D9" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- CMP a,Y
            when X"DA" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"DB" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"DC" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"DD" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- CMP a,X
            when X"DE" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- DEC a,X
            when X"DF" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";

            when X"E0" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- CPX #
            when X"E1" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- SBC (d,X)
            when X"E2" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"E3" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"E4" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- CPX d
            when X"E5" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- SBC d
            when X"E6" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- INC d
            when X"E7" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"E8" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- INX
            when X"E9" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- SBC #
            when X"EA" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- NOP
            when X"EB" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"EC" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- CPX a
            when X"ED" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- SBC a
            when X"EE" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- INC a
            when X"EF" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";

            when X"F0" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- BEQ r
            when X"F1" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- SBC (d),Y
            when X"F2" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"F3" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"F4" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"F5" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- SBC d,X
            when X"F6" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- INC d,X
            when X"F7" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"F8" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- SED
            when X"F9" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- SBC a,Y
            when X"FA" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"FB" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"FC" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"FD" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- SBC a,X
            when X"FE" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- INC a,X
            when X"FF" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";

            when others =>ctl <= B"0_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; 
         end case;
      end if;

      if cnt_r = 6 then
         case inst_r is
            when X"00" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- BRK b
            when X"01" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ORA (d,X)
            when X"02" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"03" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"04" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"05" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ORA d
            when X"06" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ASL d
            when X"07" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"08" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- PHP
            when X"09" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ORA #
            when X"0A" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ASL A
            when X"0B" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"0C" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"0D" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ORA a
            when X"0E" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ASL a
            when X"0F" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";

            when X"10" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- BPL r
            when X"11" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ORA (d),Y
            when X"12" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"13" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"14" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"15" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ORA d,X
            when X"16" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ASL d,X
            when X"17" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"18" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- CLC
            when X"19" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ORA a,Y
            when X"1A" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"1B" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"1C" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"1D" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ORA a,X
            when X"1E" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ASL a,X
            when X"1F" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";

            when X"20" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- JSR a
            when X"21" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- AND (d,X)
            when X"22" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"23" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"24" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- BIT d
            when X"25" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- AND d
            when X"26" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ROL d
            when X"27" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"28" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- PLP
            when X"29" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- AND #
            when X"2A" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ROL A
            when X"2B" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"2C" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- BIT a
            when X"2D" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- AND a
            when X"2E" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ROL a
            when X"2F" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";

            when X"30" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- BMI r
            when X"31" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- AND (d),Y
            when X"32" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"33" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"34" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"35" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- AND d,X
            when X"36" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ROL d,X
            when X"37" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"38" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- SEC
            when X"39" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- AND a,Y
            when X"3A" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"3B" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"3C" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"3D" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- AND a,X
            when X"3E" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ROL a,X
            when X"3F" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";

            when X"40" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- RTI
            when X"41" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- EOR (d,X)
            when X"42" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"43" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"44" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"45" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- EOR d
            when X"46" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LSR d
            when X"47" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"48" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- PHA
            when X"49" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- EOR #
            when X"4A" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LSR A
            when X"4B" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"4C" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- JMP a
            when X"4D" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- EOR a
            when X"4E" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LSR a
            when X"4F" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";

            when X"50" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- BVC r
            when X"51" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- EOR (d),Y
            when X"52" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"53" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"54" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"55" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- EOR d,X
            when X"56" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LSR d,X
            when X"57" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"58" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- CLI
            when X"59" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- EOR a,Y
            when X"5A" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"5B" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"5C" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"5D" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- EOR a,X
            when X"5E" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LSR a,X
            when X"5F" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";

            when X"60" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- RTS
            when X"61" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ADC (d,X)
            when X"62" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"63" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"64" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"65" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ADC d
            when X"66" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ROR d
            when X"67" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"68" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- PLA
            when X"69" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ADC #
            when X"6A" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ROR A
            when X"6B" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"6C" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- JMP (a)
            when X"6D" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ADC a
            when X"6E" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ROR a
            when X"6F" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";

            when X"70" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- BVS r
            when X"71" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ADC (d),Y
            when X"72" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"73" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"74" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"75" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ADC d,X
            when X"76" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ROR d,X
            when X"77" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"78" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- SEI
            when X"79" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ADC a,Y
            when X"7A" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"7B" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"7C" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"7D" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ADC a,X
            when X"7E" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ROR a,X
            when X"7F" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";

            when X"80" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"81" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- STA (d,X)
            when X"82" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"83" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"84" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- STY
            when X"85" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- STA d
            when X"86" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- STX d
            when X"87" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"88" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- DEY
            when X"89" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"8A" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- TXA
            when X"8B" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; 
            when X"8C" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- STY a
            when X"8D" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- STA a
            when X"8E" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- STX a
            when X"8F" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";

            when X"90" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- BCC r
            when X"91" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- STA (d),Y
            when X"92" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"93" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"94" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- STY d,X
            when X"95" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- STA d,X
            when X"96" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- STX d,Y
            when X"97" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"98" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- TYA
            when X"99" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- STA a,Y
            when X"9A" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- TXS
            when X"9B" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"9C" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"9D" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- STA a,X
            when X"9E" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"9F" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";

            when X"A0" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LDY #
            when X"A1" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LDA (d,X)
            when X"A2" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LDX #
            when X"A3" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"A4" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LDY d
            when X"A5" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LDA d
            when X"A6" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LDX d
            when X"A7" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"A8" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- TAY
            when X"A9" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LDA #
            when X"AA" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- TAX
            when X"AB" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"AC" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LDY a
            when X"AD" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LDA a
            when X"AE" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LDX a
            when X"AF" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";

            when X"B0" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- BCS r
            when X"B1" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LDA (d),Y
            when X"B2" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"B3" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"B4" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LDY d,X
            when X"B5" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LDA d,X
            when X"B6" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LDX d,Y
            when X"B7" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"B8" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- CLV
            when X"B9" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LDA a,Y
            when X"BA" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- TSX
            when X"BB" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"BC" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LDY a,X
            when X"BD" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LDA a,X
            when X"BE" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LDX a,Y
            when X"BF" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";

            when X"C0" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- CPY #
            when X"C1" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- CMP (d,X)
            when X"C2" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"C3" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"C4" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- CPY d
            when X"C5" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- CMP d
            when X"C6" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- DEC d
            when X"C7" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"C8" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- INY
            when X"C9" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- CMP #
            when X"CA" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- DEX
            when X"CB" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"CC" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- CPY a
            when X"CD" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- CMP a
            when X"CE" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- DEC a
            when X"CF" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";

            when X"D0" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- BNE r
            when X"D1" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- CMP (d),Y
            when X"D2" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"D3" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"D4" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"D5" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- CMP d,X
            when X"D6" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- DEC d,X
            when X"D7" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"D8" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- CLD
            when X"D9" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- CMP a,Y
            when X"DA" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"DB" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"DC" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"DD" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- CMP a,X
            when X"DE" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- DEC a,X
            when X"DF" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";

            when X"E0" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- CPX #
            when X"E1" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- SBC (d,X)
            when X"E2" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"E3" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"E4" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- CPX d
            when X"E5" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- SBC d
            when X"E6" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- INC d
            when X"E7" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"E8" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- INX
            when X"E9" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- SBC #
            when X"EA" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- NOP
            when X"EB" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"EC" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- CPX a
            when X"ED" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- SBC a
            when X"EE" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- INC a
            when X"EF" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";

            when X"F0" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- BEQ r
            when X"F1" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- SBC (d),Y
            when X"F2" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"F3" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"F4" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"F5" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- SBC d,X
            when X"F6" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- INC d,X
            when X"F7" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"F8" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- SED
            when X"F9" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- SBC a,Y
            when X"FA" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"FB" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"FC" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"FD" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- SBC a,X
            when X"FE" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- INC a,X
            when X"FF" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";

            when others =>ctl <= B"0_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; 
         end case;
      end if;

      if cnt_r = 7 then
         case inst_r is
            when X"00" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- BRK b
            when X"01" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ORA (d,X)
            when X"02" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"03" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"04" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"05" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ORA d
            when X"06" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ASL d
            when X"07" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"08" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- PHP
            when X"09" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ORA #
            when X"0A" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ASL A
            when X"0B" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"0C" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"0D" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ORA a
            when X"0E" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ASL a
            when X"0F" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";

            when X"10" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- BPL r
            when X"11" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ORA (d),Y
            when X"12" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"13" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"14" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"15" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ORA d,X
            when X"16" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ASL d,X
            when X"17" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"18" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- CLC
            when X"19" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ORA a,Y
            when X"1A" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"1B" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"1C" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"1D" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ORA a,X
            when X"1E" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ASL a,X
            when X"1F" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";

            when X"20" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- JSR a
            when X"21" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- AND (d,X)
            when X"22" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"23" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"24" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- BIT d
            when X"25" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- AND d
            when X"26" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ROL d
            when X"27" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"28" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- PLP
            when X"29" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- AND #
            when X"2A" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ROL A
            when X"2B" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"2C" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- BIT a
            when X"2D" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- AND a
            when X"2E" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ROL a
            when X"2F" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";

            when X"30" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- BMI r
            when X"31" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- AND (d),Y
            when X"32" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"33" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"34" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"35" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- AND d,X
            when X"36" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ROL d,X
            when X"37" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"38" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- SEC
            when X"39" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- AND a,Y
            when X"3A" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"3B" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"3C" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"3D" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- AND a,X
            when X"3E" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ROL a,X
            when X"3F" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";

            when X"40" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- RTI
            when X"41" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- EOR (d,X)
            when X"42" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"43" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"44" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"45" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- EOR d
            when X"46" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LSR d
            when X"47" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"48" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- PHA
            when X"49" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- EOR #
            when X"4A" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LSR A
            when X"4B" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"4C" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- JMP a
            when X"4D" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- EOR a
            when X"4E" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LSR a
            when X"4F" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";

            when X"50" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- BVC r
            when X"51" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- EOR (d),Y
            when X"52" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"53" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"54" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"55" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- EOR d,X
            when X"56" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LSR d,X
            when X"57" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"58" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- CLI
            when X"59" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- EOR a,Y
            when X"5A" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"5B" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"5C" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"5D" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- EOR a,X
            when X"5E" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LSR a,X
            when X"5F" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";

            when X"60" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- RTS
            when X"61" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ADC (d,X)
            when X"62" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"63" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"64" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"65" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ADC d
            when X"66" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ROR d
            when X"67" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"68" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- PLA
            when X"69" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ADC #
            when X"6A" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ROR A
            when X"6B" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"6C" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- JMP (a)
            when X"6D" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ADC a
            when X"6E" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ROR a
            when X"6F" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";

            when X"70" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- BVS r
            when X"71" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ADC (d),Y
            when X"72" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"73" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"74" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"75" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ADC d,X
            when X"76" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ROR d,X
            when X"77" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"78" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- SEI
            when X"79" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ADC a,Y
            when X"7A" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"7B" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"7C" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"7D" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ADC a,X
            when X"7E" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- ROR a,X
            when X"7F" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";

            when X"80" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"81" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- STA (d,X)
            when X"82" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"83" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"84" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- STY
            when X"85" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- STA d
            when X"86" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- STX d
            when X"87" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"88" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- DEY
            when X"89" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"8A" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- TXA
            when X"8B" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; 
            when X"8C" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- STY a
            when X"8D" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- STA a
            when X"8E" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- STX a
            when X"8F" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";

            when X"90" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- BCC r
            when X"91" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- STA (d),Y
            when X"92" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"93" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"94" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- STY d,X
            when X"95" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- STA d,X
            when X"96" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- STX d,Y
            when X"97" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"98" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- TYA
            when X"99" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- STA a,Y
            when X"9A" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- TXS
            when X"9B" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"9C" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"9D" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- STA a,X
            when X"9E" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"9F" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";

            when X"A0" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LDY #
            when X"A1" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LDA (d,X)
            when X"A2" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LDX #
            when X"A3" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"A4" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LDY d
            when X"A5" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LDA d
            when X"A6" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LDX d
            when X"A7" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"A8" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- TAY
            when X"A9" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LDA #
            when X"AA" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- TAX
            when X"AB" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"AC" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LDY a
            when X"AD" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LDA a
            when X"AE" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LDX a
            when X"AF" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";

            when X"B0" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- BCS r
            when X"B1" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LDA (d),Y
            when X"B2" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"B3" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"B4" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LDY d,X
            when X"B5" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LDA d,X
            when X"B6" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LDX d,Y
            when X"B7" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"B8" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- CLV
            when X"B9" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LDA a,Y
            when X"BA" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- TSX
            when X"BB" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"BC" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LDY a,X
            when X"BD" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LDA a,X
            when X"BE" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- LDX a,Y
            when X"BF" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";

            when X"C0" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- CPY #
            when X"C1" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- CMP (d,X)
            when X"C2" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"C3" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"C4" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- CPY d
            when X"C5" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- CMP d
            when X"C6" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- DEC d
            when X"C7" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"C8" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- INY
            when X"C9" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- CMP #
            when X"CA" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- DEX
            when X"CB" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"CC" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- CPY a
            when X"CD" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- CMP a
            when X"CE" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- DEC a
            when X"CF" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";

            when X"D0" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- BNE r
            when X"D1" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- CMP (d),Y
            when X"D2" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"D3" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"D4" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"D5" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- CMP d,X
            when X"D6" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- DEC d,X
            when X"D7" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"D8" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- CLD
            when X"D9" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- CMP a,Y
            when X"DA" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"DB" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"DC" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"DD" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- CMP a,X
            when X"DE" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- DEC a,X
            when X"DF" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";

            when X"E0" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- CPX #
            when X"E1" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- SBC (d,X)
            when X"E2" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"E3" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"E4" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- CPX d
            when X"E5" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- SBC d
            when X"E6" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- INC d
            when X"E7" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"E8" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- INX
            when X"E9" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- SBC #
            when X"EA" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- NOP
            when X"EB" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"EC" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- CPX a
            when X"ED" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- SBC a
            when X"EE" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- INC a
            when X"EF" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";

            when X"F0" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- BEQ r
            when X"F1" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- SBC (d),Y
            when X"F2" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"F3" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"F4" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"F5" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- SBC d,X
            when X"F6" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- INC d,X
            when X"F7" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"F8" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- SED
            when X"F9" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- SBC a,Y
            when X"FA" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"FB" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"FC" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";
            when X"FD" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- SBC a,X
            when X"FE" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; -- INC a,X
            when X"FF" => ctl <= B"1_0_0_0_0000_00_00_00_0_00_0000_0_0_0";

            when others =>ctl <= B"0_0_0_0_0000_00_00_00_0_00_0000_0_0_0"; 
         end case;
      end if;

   end process;

end architecture Structural;

